module AD_Table(Data_In,BCD_Out,Table_CLK);

input Table_CLK;
input [11:0]Data_In;
output [11:0]BCD_Out;

reg [11:0]BCD_Out;


always@(posedge Table_CLK)
begin
	case(Data_In)
		12'd0:BCD_Out <= 12'b000000000000;
		12'd1:BCD_Out <= 12'b000000000000;
		12'd2:BCD_Out <= 12'b000000000000;
		12'd3:BCD_Out <= 12'b000000000000;
		12'd4:BCD_Out <= 12'b000000000000;
		12'd5:BCD_Out <= 12'b000000000000;
		12'd6:BCD_Out <= 12'b000000000000;
		12'd7:BCD_Out <= 12'b000000000000;
		12'd8:BCD_Out <= 12'b000000000000;
		12'd9:BCD_Out <= 12'b000000000001;
		12'd10:BCD_Out <= 12'b000000000001;
		12'd11:BCD_Out <= 12'b000000000001;
		12'd12:BCD_Out <= 12'b000000000001;
		12'd13:BCD_Out <= 12'b000000000001;
		12'd14:BCD_Out <= 12'b000000000001;
		12'd15:BCD_Out <= 12'b000000000001;
		12'd16:BCD_Out <= 12'b000000000001;
		12'd17:BCD_Out <= 12'b000000000001;
		12'd18:BCD_Out <= 12'b000000000001;
		12'd19:BCD_Out <= 12'b000000000001;
		12'd20:BCD_Out <= 12'b000000000001;
		12'd21:BCD_Out <= 12'b000000000001;
		12'd22:BCD_Out <= 12'b000000000001;
		12'd23:BCD_Out <= 12'b000000000001;
		12'd24:BCD_Out <= 12'b000000000001;
		12'd25:BCD_Out <= 12'b000000000010;
		12'd26:BCD_Out <= 12'b000000000010;
		12'd27:BCD_Out <= 12'b000000000010;
		12'd28:BCD_Out <= 12'b000000000010;
		12'd29:BCD_Out <= 12'b000000000010;
		12'd30:BCD_Out <= 12'b000000000010;
		12'd31:BCD_Out <= 12'b000000000010;
		12'd32:BCD_Out <= 12'b000000000010;
		12'd33:BCD_Out <= 12'b000000000010;
		12'd34:BCD_Out <= 12'b000000000010;
		12'd35:BCD_Out <= 12'b000000000010;
		12'd36:BCD_Out <= 12'b000000000010;
		12'd37:BCD_Out <= 12'b000000000010;
		12'd38:BCD_Out <= 12'b000000000010;
		12'd39:BCD_Out <= 12'b000000000010;
		12'd40:BCD_Out <= 12'b000000000010;
		12'd41:BCD_Out <= 12'b000000000011;
		12'd42:BCD_Out <= 12'b000000000011;
		12'd43:BCD_Out <= 12'b000000000011;
		12'd44:BCD_Out <= 12'b000000000011;
		12'd45:BCD_Out <= 12'b000000000011;
		12'd46:BCD_Out <= 12'b000000000011;
		12'd47:BCD_Out <= 12'b000000000011;
		12'd48:BCD_Out <= 12'b000000000011;
		12'd49:BCD_Out <= 12'b000000000011;
		12'd50:BCD_Out <= 12'b000000000011;
		12'd51:BCD_Out <= 12'b000000000011;
		12'd52:BCD_Out <= 12'b000000000011;
		12'd53:BCD_Out <= 12'b000000000011;
		12'd54:BCD_Out <= 12'b000000000011;
		12'd55:BCD_Out <= 12'b000000000011;
		12'd56:BCD_Out <= 12'b000000000011;
		12'd57:BCD_Out <= 12'b000000000011;
		12'd58:BCD_Out <= 12'b000000000100;
		12'd59:BCD_Out <= 12'b000000000100;
		12'd60:BCD_Out <= 12'b000000000100;
		12'd61:BCD_Out <= 12'b000000000100;
		12'd62:BCD_Out <= 12'b000000000100;
		12'd63:BCD_Out <= 12'b000000000100;
		12'd64:BCD_Out <= 12'b000000000100;
		12'd65:BCD_Out <= 12'b000000000100;
		12'd66:BCD_Out <= 12'b000000000100;
		12'd67:BCD_Out <= 12'b000000000100;
		12'd68:BCD_Out <= 12'b000000000100;
		12'd69:BCD_Out <= 12'b000000000100;
		12'd70:BCD_Out <= 12'b000000000100;
		12'd71:BCD_Out <= 12'b000000000100;
		12'd72:BCD_Out <= 12'b000000000100;
		12'd73:BCD_Out <= 12'b000000000100;
		12'd74:BCD_Out <= 12'b000000000101;
		12'd75:BCD_Out <= 12'b000000000101;
		12'd76:BCD_Out <= 12'b000000000101;
		12'd77:BCD_Out <= 12'b000000000101;
		12'd78:BCD_Out <= 12'b000000000101;
		12'd79:BCD_Out <= 12'b000000000101;
		12'd80:BCD_Out <= 12'b000000000101;
		12'd81:BCD_Out <= 12'b000000000101;
		12'd82:BCD_Out <= 12'b000000000101;
		12'd83:BCD_Out <= 12'b000000000101;
		12'd84:BCD_Out <= 12'b000000000101;
		12'd85:BCD_Out <= 12'b000000000101;
		12'd86:BCD_Out <= 12'b000000000101;
		12'd87:BCD_Out <= 12'b000000000101;
		12'd88:BCD_Out <= 12'b000000000101;
		12'd89:BCD_Out <= 12'b000000000101;
		12'd90:BCD_Out <= 12'b000000000101;
		12'd91:BCD_Out <= 12'b000000000110;
		12'd92:BCD_Out <= 12'b000000000110;
		12'd93:BCD_Out <= 12'b000000000110;
		12'd94:BCD_Out <= 12'b000000000110;
		12'd95:BCD_Out <= 12'b000000000110;
		12'd96:BCD_Out <= 12'b000000000110;
		12'd97:BCD_Out <= 12'b000000000110;
		12'd98:BCD_Out <= 12'b000000000110;
		12'd99:BCD_Out <= 12'b000000000110;
		12'd100:BCD_Out <= 12'b000000000110;
		12'd101:BCD_Out <= 12'b000000000110;
		12'd102:BCD_Out <= 12'b000000000110;
		12'd103:BCD_Out <= 12'b000000000110;
		12'd104:BCD_Out <= 12'b000000000110;
		12'd105:BCD_Out <= 12'b000000000110;
		12'd106:BCD_Out <= 12'b000000000110;
		12'd107:BCD_Out <= 12'b000000000111;
		12'd108:BCD_Out <= 12'b000000000111;
		12'd109:BCD_Out <= 12'b000000000111;
		12'd110:BCD_Out <= 12'b000000000111;
		12'd111:BCD_Out <= 12'b000000000111;
		12'd112:BCD_Out <= 12'b000000000111;
		12'd113:BCD_Out <= 12'b000000000111;
		12'd114:BCD_Out <= 12'b000000000111;
		12'd115:BCD_Out <= 12'b000000000111;
		12'd116:BCD_Out <= 12'b000000000111;
		12'd117:BCD_Out <= 12'b000000000111;
		12'd118:BCD_Out <= 12'b000000000111;
		12'd119:BCD_Out <= 12'b000000000111;
		12'd120:BCD_Out <= 12'b000000000111;
		12'd121:BCD_Out <= 12'b000000000111;
		12'd122:BCD_Out <= 12'b000000000111;
		12'd123:BCD_Out <= 12'b000000001000;
		12'd124:BCD_Out <= 12'b000000001000;
		12'd125:BCD_Out <= 12'b000000001000;
		12'd126:BCD_Out <= 12'b000000001000;
		12'd127:BCD_Out <= 12'b000000001000;
		12'd128:BCD_Out <= 12'b000000001000;
		12'd129:BCD_Out <= 12'b000000001000;
		12'd130:BCD_Out <= 12'b000000001000;
		12'd131:BCD_Out <= 12'b000000001000;
		12'd132:BCD_Out <= 12'b000000001000;
		12'd133:BCD_Out <= 12'b000000001000;
		12'd134:BCD_Out <= 12'b000000001000;
		12'd135:BCD_Out <= 12'b000000001000;
		12'd136:BCD_Out <= 12'b000000001000;
		12'd137:BCD_Out <= 12'b000000001000;
		12'd138:BCD_Out <= 12'b000000001000;
		12'd139:BCD_Out <= 12'b000000001000;
		12'd140:BCD_Out <= 12'b000000001001;
		12'd141:BCD_Out <= 12'b000000001001;
		12'd142:BCD_Out <= 12'b000000001001;
		12'd143:BCD_Out <= 12'b000000001001;
		12'd144:BCD_Out <= 12'b000000001001;
		12'd145:BCD_Out <= 12'b000000001001;
		12'd146:BCD_Out <= 12'b000000001001;
		12'd147:BCD_Out <= 12'b000000001001;
		12'd148:BCD_Out <= 12'b000000001001;
		12'd149:BCD_Out <= 12'b000000001001;
		12'd150:BCD_Out <= 12'b000000001001;
		12'd151:BCD_Out <= 12'b000000001001;
		12'd152:BCD_Out <= 12'b000000001001;
		12'd153:BCD_Out <= 12'b000000001001;
		12'd154:BCD_Out <= 12'b000000001001;
		12'd155:BCD_Out <= 12'b000000001001;
		12'd156:BCD_Out <= 12'b000000010000;
		12'd157:BCD_Out <= 12'b000000010000;
		12'd158:BCD_Out <= 12'b000000010000;
		12'd159:BCD_Out <= 12'b000000010000;
		12'd160:BCD_Out <= 12'b000000010000;
		12'd161:BCD_Out <= 12'b000000010000;
		12'd162:BCD_Out <= 12'b000000010000;
		12'd163:BCD_Out <= 12'b000000010000;
		12'd164:BCD_Out <= 12'b000000010000;
		12'd165:BCD_Out <= 12'b000000010000;
		12'd166:BCD_Out <= 12'b000000010000;
		12'd167:BCD_Out <= 12'b000000010000;
		12'd168:BCD_Out <= 12'b000000010000;
		12'd169:BCD_Out <= 12'b000000010000;
		12'd170:BCD_Out <= 12'b000000010000;
		12'd171:BCD_Out <= 12'b000000010000;
		12'd172:BCD_Out <= 12'b000000010001;
		12'd173:BCD_Out <= 12'b000000010001;
		12'd174:BCD_Out <= 12'b000000010001;
		12'd175:BCD_Out <= 12'b000000010001;
		12'd176:BCD_Out <= 12'b000000010001;
		12'd177:BCD_Out <= 12'b000000010001;
		12'd178:BCD_Out <= 12'b000000010001;
		12'd179:BCD_Out <= 12'b000000010001;
		12'd180:BCD_Out <= 12'b000000010001;
		12'd181:BCD_Out <= 12'b000000010001;
		12'd182:BCD_Out <= 12'b000000010001;
		12'd183:BCD_Out <= 12'b000000010001;
		12'd184:BCD_Out <= 12'b000000010001;
		12'd185:BCD_Out <= 12'b000000010001;
		12'd186:BCD_Out <= 12'b000000010001;
		12'd187:BCD_Out <= 12'b000000010001;
		12'd188:BCD_Out <= 12'b000000010001;
		12'd189:BCD_Out <= 12'b000000010010;
		12'd190:BCD_Out <= 12'b000000010010;
		12'd191:BCD_Out <= 12'b000000010010;
		12'd192:BCD_Out <= 12'b000000010010;
		12'd193:BCD_Out <= 12'b000000010010;
		12'd194:BCD_Out <= 12'b000000010010;
		12'd195:BCD_Out <= 12'b000000010010;
		12'd196:BCD_Out <= 12'b000000010010;
		12'd197:BCD_Out <= 12'b000000010010;
		12'd198:BCD_Out <= 12'b000000010010;
		12'd199:BCD_Out <= 12'b000000010010;
		12'd200:BCD_Out <= 12'b000000010010;
		12'd201:BCD_Out <= 12'b000000010010;
		12'd202:BCD_Out <= 12'b000000010010;
		12'd203:BCD_Out <= 12'b000000010010;
		12'd204:BCD_Out <= 12'b000000010010;
		12'd205:BCD_Out <= 12'b000000010011;
		12'd206:BCD_Out <= 12'b000000010011;
		12'd207:BCD_Out <= 12'b000000010011;
		12'd208:BCD_Out <= 12'b000000010011;
		12'd209:BCD_Out <= 12'b000000010011;
		12'd210:BCD_Out <= 12'b000000010011;
		12'd211:BCD_Out <= 12'b000000010011;
		12'd212:BCD_Out <= 12'b000000010011;
		12'd213:BCD_Out <= 12'b000000010011;
		12'd214:BCD_Out <= 12'b000000010011;
		12'd215:BCD_Out <= 12'b000000010011;
		12'd216:BCD_Out <= 12'b000000010011;
		12'd217:BCD_Out <= 12'b000000010011;
		12'd218:BCD_Out <= 12'b000000010011;
		12'd219:BCD_Out <= 12'b000000010011;
		12'd220:BCD_Out <= 12'b000000010011;
		12'd221:BCD_Out <= 12'b000000010011;
		12'd222:BCD_Out <= 12'b000000010100;
		12'd223:BCD_Out <= 12'b000000010100;
		12'd224:BCD_Out <= 12'b000000010100;
		12'd225:BCD_Out <= 12'b000000010100;
		12'd226:BCD_Out <= 12'b000000010100;
		12'd227:BCD_Out <= 12'b000000010100;
		12'd228:BCD_Out <= 12'b000000010100;
		12'd229:BCD_Out <= 12'b000000010100;
		12'd230:BCD_Out <= 12'b000000010100;
		12'd231:BCD_Out <= 12'b000000010100;
		12'd232:BCD_Out <= 12'b000000010100;
		12'd233:BCD_Out <= 12'b000000010100;
		12'd234:BCD_Out <= 12'b000000010100;
		12'd235:BCD_Out <= 12'b000000010100;
		12'd236:BCD_Out <= 12'b000000010100;
		12'd237:BCD_Out <= 12'b000000010100;
		12'd238:BCD_Out <= 12'b000000010101;
		12'd239:BCD_Out <= 12'b000000010101;
		12'd240:BCD_Out <= 12'b000000010101;
		12'd241:BCD_Out <= 12'b000000010101;
		12'd242:BCD_Out <= 12'b000000010101;
		12'd243:BCD_Out <= 12'b000000010101;
		12'd244:BCD_Out <= 12'b000000010101;
		12'd245:BCD_Out <= 12'b000000010101;
		12'd246:BCD_Out <= 12'b000000010101;
		12'd247:BCD_Out <= 12'b000000010101;
		12'd248:BCD_Out <= 12'b000000010101;
		12'd249:BCD_Out <= 12'b000000010101;
		12'd250:BCD_Out <= 12'b000000010101;
		12'd251:BCD_Out <= 12'b000000010101;
		12'd252:BCD_Out <= 12'b000000010101;
		12'd253:BCD_Out <= 12'b000000010101;
		12'd254:BCD_Out <= 12'b000000010110;
		12'd255:BCD_Out <= 12'b000000010110;
		12'd256:BCD_Out <= 12'b000000010110;
		12'd257:BCD_Out <= 12'b000000010110;
		12'd258:BCD_Out <= 12'b000000010110;
		12'd259:BCD_Out <= 12'b000000010110;
		12'd260:BCD_Out <= 12'b000000010110;
		12'd261:BCD_Out <= 12'b000000010110;
		12'd262:BCD_Out <= 12'b000000010110;
		12'd263:BCD_Out <= 12'b000000010110;
		12'd264:BCD_Out <= 12'b000000010110;
		12'd265:BCD_Out <= 12'b000000010110;
		12'd266:BCD_Out <= 12'b000000010110;
		12'd267:BCD_Out <= 12'b000000010110;
		12'd268:BCD_Out <= 12'b000000010110;
		12'd269:BCD_Out <= 12'b000000010110;
		12'd270:BCD_Out <= 12'b000000010110;
		12'd271:BCD_Out <= 12'b000000010111;
		12'd272:BCD_Out <= 12'b000000010111;
		12'd273:BCD_Out <= 12'b000000010111;
		12'd274:BCD_Out <= 12'b000000010111;
		12'd275:BCD_Out <= 12'b000000010111;
		12'd276:BCD_Out <= 12'b000000010111;
		12'd277:BCD_Out <= 12'b000000010111;
		12'd278:BCD_Out <= 12'b000000010111;
		12'd279:BCD_Out <= 12'b000000010111;
		12'd280:BCD_Out <= 12'b000000010111;
		12'd281:BCD_Out <= 12'b000000010111;
		12'd282:BCD_Out <= 12'b000000010111;
		12'd283:BCD_Out <= 12'b000000010111;
		12'd284:BCD_Out <= 12'b000000010111;
		12'd285:BCD_Out <= 12'b000000010111;
		12'd286:BCD_Out <= 12'b000000010111;
		12'd287:BCD_Out <= 12'b000000011000;
		12'd288:BCD_Out <= 12'b000000011000;
		12'd289:BCD_Out <= 12'b000000011000;
		12'd290:BCD_Out <= 12'b000000011000;
		12'd291:BCD_Out <= 12'b000000011000;
		12'd292:BCD_Out <= 12'b000000011000;
		12'd293:BCD_Out <= 12'b000000011000;
		12'd294:BCD_Out <= 12'b000000011000;
		12'd295:BCD_Out <= 12'b000000011000;
		12'd296:BCD_Out <= 12'b000000011000;
		12'd297:BCD_Out <= 12'b000000011000;
		12'd298:BCD_Out <= 12'b000000011000;
		12'd299:BCD_Out <= 12'b000000011000;
		12'd300:BCD_Out <= 12'b000000011000;
		12'd301:BCD_Out <= 12'b000000011000;
		12'd302:BCD_Out <= 12'b000000011000;
		12'd303:BCD_Out <= 12'b000000011000;
		12'd304:BCD_Out <= 12'b000000011001;
		12'd305:BCD_Out <= 12'b000000011001;
		12'd306:BCD_Out <= 12'b000000011001;
		12'd307:BCD_Out <= 12'b000000011001;
		12'd308:BCD_Out <= 12'b000000011001;
		12'd309:BCD_Out <= 12'b000000011001;
		12'd310:BCD_Out <= 12'b000000011001;
		12'd311:BCD_Out <= 12'b000000011001;
		12'd312:BCD_Out <= 12'b000000011001;
		12'd313:BCD_Out <= 12'b000000011001;
		12'd314:BCD_Out <= 12'b000000011001;
		12'd315:BCD_Out <= 12'b000000011001;
		12'd316:BCD_Out <= 12'b000000011001;
		12'd317:BCD_Out <= 12'b000000011001;
		12'd318:BCD_Out <= 12'b000000011001;
		12'd319:BCD_Out <= 12'b000000011001;
		12'd320:BCD_Out <= 12'b000000100000;
		12'd321:BCD_Out <= 12'b000000100000;
		12'd322:BCD_Out <= 12'b000000100000;
		12'd323:BCD_Out <= 12'b000000100000;
		12'd324:BCD_Out <= 12'b000000100000;
		12'd325:BCD_Out <= 12'b000000100000;
		12'd326:BCD_Out <= 12'b000000100000;
		12'd327:BCD_Out <= 12'b000000100000;
		12'd328:BCD_Out <= 12'b000000100000;
		12'd329:BCD_Out <= 12'b000000100000;
		12'd330:BCD_Out <= 12'b000000100000;
		12'd331:BCD_Out <= 12'b000000100000;
		12'd332:BCD_Out <= 12'b000000100000;
		12'd333:BCD_Out <= 12'b000000100000;
		12'd334:BCD_Out <= 12'b000000100000;
		12'd335:BCD_Out <= 12'b000000100000;
		12'd336:BCD_Out <= 12'b000000100001;
		12'd337:BCD_Out <= 12'b000000100001;
		12'd338:BCD_Out <= 12'b000000100001;
		12'd339:BCD_Out <= 12'b000000100001;
		12'd340:BCD_Out <= 12'b000000100001;
		12'd341:BCD_Out <= 12'b000000100001;
		12'd342:BCD_Out <= 12'b000000100001;
		12'd343:BCD_Out <= 12'b000000100001;
		12'd344:BCD_Out <= 12'b000000100001;
		12'd345:BCD_Out <= 12'b000000100001;
		12'd346:BCD_Out <= 12'b000000100001;
		12'd347:BCD_Out <= 12'b000000100001;
		12'd348:BCD_Out <= 12'b000000100001;
		12'd349:BCD_Out <= 12'b000000100001;
		12'd350:BCD_Out <= 12'b000000100001;
		12'd351:BCD_Out <= 12'b000000100001;
		12'd352:BCD_Out <= 12'b000000100001;
		12'd353:BCD_Out <= 12'b000000100010;
		12'd354:BCD_Out <= 12'b000000100010;
		12'd355:BCD_Out <= 12'b000000100010;
		12'd356:BCD_Out <= 12'b000000100010;
		12'd357:BCD_Out <= 12'b000000100010;
		12'd358:BCD_Out <= 12'b000000100010;
		12'd359:BCD_Out <= 12'b000000100010;
		12'd360:BCD_Out <= 12'b000000100010;
		12'd361:BCD_Out <= 12'b000000100010;
		12'd362:BCD_Out <= 12'b000000100010;
		12'd363:BCD_Out <= 12'b000000100010;
		12'd364:BCD_Out <= 12'b000000100010;
		12'd365:BCD_Out <= 12'b000000100010;
		12'd366:BCD_Out <= 12'b000000100010;
		12'd367:BCD_Out <= 12'b000000100010;
		12'd368:BCD_Out <= 12'b000000100010;
		12'd369:BCD_Out <= 12'b000000100011;
		12'd370:BCD_Out <= 12'b000000100011;
		12'd371:BCD_Out <= 12'b000000100011;
		12'd372:BCD_Out <= 12'b000000100011;
		12'd373:BCD_Out <= 12'b000000100011;
		12'd374:BCD_Out <= 12'b000000100011;
		12'd375:BCD_Out <= 12'b000000100011;
		12'd376:BCD_Out <= 12'b000000100011;
		12'd377:BCD_Out <= 12'b000000100011;
		12'd378:BCD_Out <= 12'b000000100011;
		12'd379:BCD_Out <= 12'b000000100011;
		12'd380:BCD_Out <= 12'b000000100011;
		12'd381:BCD_Out <= 12'b000000100011;
		12'd382:BCD_Out <= 12'b000000100011;
		12'd383:BCD_Out <= 12'b000000100011;
		12'd384:BCD_Out <= 12'b000000100011;
		12'd385:BCD_Out <= 12'b000000100100;
		12'd386:BCD_Out <= 12'b000000100100;
		12'd387:BCD_Out <= 12'b000000100100;
		12'd388:BCD_Out <= 12'b000000100100;
		12'd389:BCD_Out <= 12'b000000100100;
		12'd390:BCD_Out <= 12'b000000100100;
		12'd391:BCD_Out <= 12'b000000100100;
		12'd392:BCD_Out <= 12'b000000100100;
		12'd393:BCD_Out <= 12'b000000100100;
		12'd394:BCD_Out <= 12'b000000100100;
		12'd395:BCD_Out <= 12'b000000100100;
		12'd396:BCD_Out <= 12'b000000100100;
		12'd397:BCD_Out <= 12'b000000100100;
		12'd398:BCD_Out <= 12'b000000100100;
		12'd399:BCD_Out <= 12'b000000100100;
		12'd400:BCD_Out <= 12'b000000100100;
		12'd401:BCD_Out <= 12'b000000100100;
		12'd402:BCD_Out <= 12'b000000100101;
		12'd403:BCD_Out <= 12'b000000100101;
		12'd404:BCD_Out <= 12'b000000100101;
		12'd405:BCD_Out <= 12'b000000100101;
		12'd406:BCD_Out <= 12'b000000100101;
		12'd407:BCD_Out <= 12'b000000100101;
		12'd408:BCD_Out <= 12'b000000100101;
		12'd409:BCD_Out <= 12'b000000100101;
		12'd410:BCD_Out <= 12'b000000100101;
		12'd411:BCD_Out <= 12'b000000100101;
		12'd412:BCD_Out <= 12'b000000100101;
		12'd413:BCD_Out <= 12'b000000100101;
		12'd414:BCD_Out <= 12'b000000100101;
		12'd415:BCD_Out <= 12'b000000100101;
		12'd416:BCD_Out <= 12'b000000100101;
		12'd417:BCD_Out <= 12'b000000100101;
		12'd418:BCD_Out <= 12'b000000100110;
		12'd419:BCD_Out <= 12'b000000100110;
		12'd420:BCD_Out <= 12'b000000100110;
		12'd421:BCD_Out <= 12'b000000100110;
		12'd422:BCD_Out <= 12'b000000100110;
		12'd423:BCD_Out <= 12'b000000100110;
		12'd424:BCD_Out <= 12'b000000100110;
		12'd425:BCD_Out <= 12'b000000100110;
		12'd426:BCD_Out <= 12'b000000100110;
		12'd427:BCD_Out <= 12'b000000100110;
		12'd428:BCD_Out <= 12'b000000100110;
		12'd429:BCD_Out <= 12'b000000100110;
		12'd430:BCD_Out <= 12'b000000100110;
		12'd431:BCD_Out <= 12'b000000100110;
		12'd432:BCD_Out <= 12'b000000100110;
		12'd433:BCD_Out <= 12'b000000100110;
		12'd434:BCD_Out <= 12'b000000100110;
		12'd435:BCD_Out <= 12'b000000100111;
		12'd436:BCD_Out <= 12'b000000100111;
		12'd437:BCD_Out <= 12'b000000100111;
		12'd438:BCD_Out <= 12'b000000100111;
		12'd439:BCD_Out <= 12'b000000100111;
		12'd440:BCD_Out <= 12'b000000100111;
		12'd441:BCD_Out <= 12'b000000100111;
		12'd442:BCD_Out <= 12'b000000100111;
		12'd443:BCD_Out <= 12'b000000100111;
		12'd444:BCD_Out <= 12'b000000100111;
		12'd445:BCD_Out <= 12'b000000100111;
		12'd446:BCD_Out <= 12'b000000100111;
		12'd447:BCD_Out <= 12'b000000100111;
		12'd448:BCD_Out <= 12'b000000100111;
		12'd449:BCD_Out <= 12'b000000100111;
		12'd450:BCD_Out <= 12'b000000100111;
		12'd451:BCD_Out <= 12'b000000101000;
		12'd452:BCD_Out <= 12'b000000101000;
		12'd453:BCD_Out <= 12'b000000101000;
		12'd454:BCD_Out <= 12'b000000101000;
		12'd455:BCD_Out <= 12'b000000101000;
		12'd456:BCD_Out <= 12'b000000101000;
		12'd457:BCD_Out <= 12'b000000101000;
		12'd458:BCD_Out <= 12'b000000101000;
		12'd459:BCD_Out <= 12'b000000101000;
		12'd460:BCD_Out <= 12'b000000101000;
		12'd461:BCD_Out <= 12'b000000101000;
		12'd462:BCD_Out <= 12'b000000101000;
		12'd463:BCD_Out <= 12'b000000101000;
		12'd464:BCD_Out <= 12'b000000101000;
		12'd465:BCD_Out <= 12'b000000101000;
		12'd466:BCD_Out <= 12'b000000101000;
		12'd467:BCD_Out <= 12'b000000101001;
		12'd468:BCD_Out <= 12'b000000101001;
		12'd469:BCD_Out <= 12'b000000101001;
		12'd470:BCD_Out <= 12'b000000101001;
		12'd471:BCD_Out <= 12'b000000101001;
		12'd472:BCD_Out <= 12'b000000101001;
		12'd473:BCD_Out <= 12'b000000101001;
		12'd474:BCD_Out <= 12'b000000101001;
		12'd475:BCD_Out <= 12'b000000101001;
		12'd476:BCD_Out <= 12'b000000101001;
		12'd477:BCD_Out <= 12'b000000101001;
		12'd478:BCD_Out <= 12'b000000101001;
		12'd479:BCD_Out <= 12'b000000101001;
		12'd480:BCD_Out <= 12'b000000101001;
		12'd481:BCD_Out <= 12'b000000101001;
		12'd482:BCD_Out <= 12'b000000101001;
		12'd483:BCD_Out <= 12'b000000101001;
		12'd484:BCD_Out <= 12'b000000110000;
		12'd485:BCD_Out <= 12'b000000110000;
		12'd486:BCD_Out <= 12'b000000110000;
		12'd487:BCD_Out <= 12'b000000110000;
		12'd488:BCD_Out <= 12'b000000110000;
		12'd489:BCD_Out <= 12'b000000110000;
		12'd490:BCD_Out <= 12'b000000110000;
		12'd491:BCD_Out <= 12'b000000110000;
		12'd492:BCD_Out <= 12'b000000110000;
		12'd493:BCD_Out <= 12'b000000110000;
		12'd494:BCD_Out <= 12'b000000110000;
		12'd495:BCD_Out <= 12'b000000110000;
		12'd496:BCD_Out <= 12'b000000110000;
		12'd497:BCD_Out <= 12'b000000110000;
		12'd498:BCD_Out <= 12'b000000110000;
		12'd499:BCD_Out <= 12'b000000110000;
		12'd500:BCD_Out <= 12'b000000110001;
		12'd501:BCD_Out <= 12'b000000110001;
		12'd502:BCD_Out <= 12'b000000110001;
		12'd503:BCD_Out <= 12'b000000110001;
		12'd504:BCD_Out <= 12'b000000110001;
		12'd505:BCD_Out <= 12'b000000110001;
		12'd506:BCD_Out <= 12'b000000110001;
		12'd507:BCD_Out <= 12'b000000110001;
		12'd508:BCD_Out <= 12'b000000110001;
		12'd509:BCD_Out <= 12'b000000110001;
		12'd510:BCD_Out <= 12'b000000110001;
		12'd511:BCD_Out <= 12'b000000110001;
		12'd512:BCD_Out <= 12'b000000110001;
		12'd513:BCD_Out <= 12'b000000110001;
		12'd514:BCD_Out <= 12'b000000110001;
		12'd515:BCD_Out <= 12'b000000110001;
		12'd516:BCD_Out <= 12'b000000110010;
		12'd517:BCD_Out <= 12'b000000110010;
		12'd518:BCD_Out <= 12'b000000110010;
		12'd519:BCD_Out <= 12'b000000110010;
		12'd520:BCD_Out <= 12'b000000110010;
		12'd521:BCD_Out <= 12'b000000110010;
		12'd522:BCD_Out <= 12'b000000110010;
		12'd523:BCD_Out <= 12'b000000110010;
		12'd524:BCD_Out <= 12'b000000110010;
		12'd525:BCD_Out <= 12'b000000110010;
		12'd526:BCD_Out <= 12'b000000110010;
		12'd527:BCD_Out <= 12'b000000110010;
		12'd528:BCD_Out <= 12'b000000110010;
		12'd529:BCD_Out <= 12'b000000110010;
		12'd530:BCD_Out <= 12'b000000110010;
		12'd531:BCD_Out <= 12'b000000110010;
		12'd532:BCD_Out <= 12'b000000110010;
		12'd533:BCD_Out <= 12'b000000110011;
		12'd534:BCD_Out <= 12'b000000110011;
		12'd535:BCD_Out <= 12'b000000110011;
		12'd536:BCD_Out <= 12'b000000110011;
		12'd537:BCD_Out <= 12'b000000110011;
		12'd538:BCD_Out <= 12'b000000110011;
		12'd539:BCD_Out <= 12'b000000110011;
		12'd540:BCD_Out <= 12'b000000110011;
		12'd541:BCD_Out <= 12'b000000110011;
		12'd542:BCD_Out <= 12'b000000110011;
		12'd543:BCD_Out <= 12'b000000110011;
		12'd544:BCD_Out <= 12'b000000110011;
		12'd545:BCD_Out <= 12'b000000110011;
		12'd546:BCD_Out <= 12'b000000110011;
		12'd547:BCD_Out <= 12'b000000110011;
		12'd548:BCD_Out <= 12'b000000110011;
		12'd549:BCD_Out <= 12'b000000110100;
		12'd550:BCD_Out <= 12'b000000110100;
		12'd551:BCD_Out <= 12'b000000110100;
		12'd552:BCD_Out <= 12'b000000110100;
		12'd553:BCD_Out <= 12'b000000110100;
		12'd554:BCD_Out <= 12'b000000110100;
		12'd555:BCD_Out <= 12'b000000110100;
		12'd556:BCD_Out <= 12'b000000110100;
		12'd557:BCD_Out <= 12'b000000110100;
		12'd558:BCD_Out <= 12'b000000110100;
		12'd559:BCD_Out <= 12'b000000110100;
		12'd560:BCD_Out <= 12'b000000110100;
		12'd561:BCD_Out <= 12'b000000110100;
		12'd562:BCD_Out <= 12'b000000110100;
		12'd563:BCD_Out <= 12'b000000110100;
		12'd564:BCD_Out <= 12'b000000110100;
		12'd565:BCD_Out <= 12'b000000110100;
		12'd566:BCD_Out <= 12'b000000110101;
		12'd567:BCD_Out <= 12'b000000110101;
		12'd568:BCD_Out <= 12'b000000110101;
		12'd569:BCD_Out <= 12'b000000110101;
		12'd570:BCD_Out <= 12'b000000110101;
		12'd571:BCD_Out <= 12'b000000110101;
		12'd572:BCD_Out <= 12'b000000110101;
		12'd573:BCD_Out <= 12'b000000110101;
		12'd574:BCD_Out <= 12'b000000110101;
		12'd575:BCD_Out <= 12'b000000110101;
		12'd576:BCD_Out <= 12'b000000110101;
		12'd577:BCD_Out <= 12'b000000110101;
		12'd578:BCD_Out <= 12'b000000110101;
		12'd579:BCD_Out <= 12'b000000110101;
		12'd580:BCD_Out <= 12'b000000110101;
		12'd581:BCD_Out <= 12'b000000110101;
		12'd582:BCD_Out <= 12'b000000110110;
		12'd583:BCD_Out <= 12'b000000110110;
		12'd584:BCD_Out <= 12'b000000110110;
		12'd585:BCD_Out <= 12'b000000110110;
		12'd586:BCD_Out <= 12'b000000110110;
		12'd587:BCD_Out <= 12'b000000110110;
		12'd588:BCD_Out <= 12'b000000110110;
		12'd589:BCD_Out <= 12'b000000110110;
		12'd590:BCD_Out <= 12'b000000110110;
		12'd591:BCD_Out <= 12'b000000110110;
		12'd592:BCD_Out <= 12'b000000110110;
		12'd593:BCD_Out <= 12'b000000110110;
		12'd594:BCD_Out <= 12'b000000110110;
		12'd595:BCD_Out <= 12'b000000110110;
		12'd596:BCD_Out <= 12'b000000110110;
		12'd597:BCD_Out <= 12'b000000110110;
		12'd598:BCD_Out <= 12'b000000110111;
		12'd599:BCD_Out <= 12'b000000110111;
		12'd600:BCD_Out <= 12'b000000110111;
		12'd601:BCD_Out <= 12'b000000110111;
		12'd602:BCD_Out <= 12'b000000110111;
		12'd603:BCD_Out <= 12'b000000110111;
		12'd604:BCD_Out <= 12'b000000110111;
		12'd605:BCD_Out <= 12'b000000110111;
		12'd606:BCD_Out <= 12'b000000110111;
		12'd607:BCD_Out <= 12'b000000110111;
		12'd608:BCD_Out <= 12'b000000110111;
		12'd609:BCD_Out <= 12'b000000110111;
		12'd610:BCD_Out <= 12'b000000110111;
		12'd611:BCD_Out <= 12'b000000110111;
		12'd612:BCD_Out <= 12'b000000110111;
		12'd613:BCD_Out <= 12'b000000110111;
		12'd614:BCD_Out <= 12'b000000110111;
		12'd615:BCD_Out <= 12'b000000111000;
		12'd616:BCD_Out <= 12'b000000111000;
		12'd617:BCD_Out <= 12'b000000111000;
		12'd618:BCD_Out <= 12'b000000111000;
		12'd619:BCD_Out <= 12'b000000111000;
		12'd620:BCD_Out <= 12'b000000111000;
		12'd621:BCD_Out <= 12'b000000111000;
		12'd622:BCD_Out <= 12'b000000111000;
		12'd623:BCD_Out <= 12'b000000111000;
		12'd624:BCD_Out <= 12'b000000111000;
		12'd625:BCD_Out <= 12'b000000111000;
		12'd626:BCD_Out <= 12'b000000111000;
		12'd627:BCD_Out <= 12'b000000111000;
		12'd628:BCD_Out <= 12'b000000111000;
		12'd629:BCD_Out <= 12'b000000111000;
		12'd630:BCD_Out <= 12'b000000111000;
		12'd631:BCD_Out <= 12'b000000111001;
		12'd632:BCD_Out <= 12'b000000111001;
		12'd633:BCD_Out <= 12'b000000111001;
		12'd634:BCD_Out <= 12'b000000111001;
		12'd635:BCD_Out <= 12'b000000111001;
		12'd636:BCD_Out <= 12'b000000111001;
		12'd637:BCD_Out <= 12'b000000111001;
		12'd638:BCD_Out <= 12'b000000111001;
		12'd639:BCD_Out <= 12'b000000111001;
		12'd640:BCD_Out <= 12'b000000111001;
		12'd641:BCD_Out <= 12'b000000111001;
		12'd642:BCD_Out <= 12'b000000111001;
		12'd643:BCD_Out <= 12'b000000111001;
		12'd644:BCD_Out <= 12'b000000111001;
		12'd645:BCD_Out <= 12'b000000111001;
		12'd646:BCD_Out <= 12'b000000111001;
		12'd647:BCD_Out <= 12'b000000111001;
		12'd648:BCD_Out <= 12'b000001000000;
		12'd649:BCD_Out <= 12'b000001000000;
		12'd650:BCD_Out <= 12'b000001000000;
		12'd651:BCD_Out <= 12'b000001000000;
		12'd652:BCD_Out <= 12'b000001000000;
		12'd653:BCD_Out <= 12'b000001000000;
		12'd654:BCD_Out <= 12'b000001000000;
		12'd655:BCD_Out <= 12'b000001000000;
		12'd656:BCD_Out <= 12'b000001000000;
		12'd657:BCD_Out <= 12'b000001000000;
		12'd658:BCD_Out <= 12'b000001000000;
		12'd659:BCD_Out <= 12'b000001000000;
		12'd660:BCD_Out <= 12'b000001000000;
		12'd661:BCD_Out <= 12'b000001000000;
		12'd662:BCD_Out <= 12'b000001000000;
		12'd663:BCD_Out <= 12'b000001000000;
		12'd664:BCD_Out <= 12'b000001000001;
		12'd665:BCD_Out <= 12'b000001000001;
		12'd666:BCD_Out <= 12'b000001000001;
		12'd667:BCD_Out <= 12'b000001000001;
		12'd668:BCD_Out <= 12'b000001000001;
		12'd669:BCD_Out <= 12'b000001000001;
		12'd670:BCD_Out <= 12'b000001000001;
		12'd671:BCD_Out <= 12'b000001000001;
		12'd672:BCD_Out <= 12'b000001000001;
		12'd673:BCD_Out <= 12'b000001000001;
		12'd674:BCD_Out <= 12'b000001000001;
		12'd675:BCD_Out <= 12'b000001000001;
		12'd676:BCD_Out <= 12'b000001000001;
		12'd677:BCD_Out <= 12'b000001000001;
		12'd678:BCD_Out <= 12'b000001000001;
		12'd679:BCD_Out <= 12'b000001000001;
		12'd680:BCD_Out <= 12'b000001000010;
		12'd681:BCD_Out <= 12'b000001000010;
		12'd682:BCD_Out <= 12'b000001000010;
		12'd683:BCD_Out <= 12'b000001000010;
		12'd684:BCD_Out <= 12'b000001000010;
		12'd685:BCD_Out <= 12'b000001000010;
		12'd686:BCD_Out <= 12'b000001000010;
		12'd687:BCD_Out <= 12'b000001000010;
		12'd688:BCD_Out <= 12'b000001000010;
		12'd689:BCD_Out <= 12'b000001000010;
		12'd690:BCD_Out <= 12'b000001000010;
		12'd691:BCD_Out <= 12'b000001000010;
		12'd692:BCD_Out <= 12'b000001000010;
		12'd693:BCD_Out <= 12'b000001000010;
		12'd694:BCD_Out <= 12'b000001000010;
		12'd695:BCD_Out <= 12'b000001000010;
		12'd696:BCD_Out <= 12'b000001000010;
		12'd697:BCD_Out <= 12'b000001000011;
		12'd698:BCD_Out <= 12'b000001000011;
		12'd699:BCD_Out <= 12'b000001000011;
		12'd700:BCD_Out <= 12'b000001000011;
		12'd701:BCD_Out <= 12'b000001000011;
		12'd702:BCD_Out <= 12'b000001000011;
		12'd703:BCD_Out <= 12'b000001000011;
		12'd704:BCD_Out <= 12'b000001000011;
		12'd705:BCD_Out <= 12'b000001000011;
		12'd706:BCD_Out <= 12'b000001000011;
		12'd707:BCD_Out <= 12'b000001000011;
		12'd708:BCD_Out <= 12'b000001000011;
		12'd709:BCD_Out <= 12'b000001000011;
		12'd710:BCD_Out <= 12'b000001000011;
		12'd711:BCD_Out <= 12'b000001000011;
		12'd712:BCD_Out <= 12'b000001000011;
		12'd713:BCD_Out <= 12'b000001000100;
		12'd714:BCD_Out <= 12'b000001000100;
		12'd715:BCD_Out <= 12'b000001000100;
		12'd716:BCD_Out <= 12'b000001000100;
		12'd717:BCD_Out <= 12'b000001000100;
		12'd718:BCD_Out <= 12'b000001000100;
		12'd719:BCD_Out <= 12'b000001000100;
		12'd720:BCD_Out <= 12'b000001000100;
		12'd721:BCD_Out <= 12'b000001000100;
		12'd722:BCD_Out <= 12'b000001000100;
		12'd723:BCD_Out <= 12'b000001000100;
		12'd724:BCD_Out <= 12'b000001000100;
		12'd725:BCD_Out <= 12'b000001000100;
		12'd726:BCD_Out <= 12'b000001000100;
		12'd727:BCD_Out <= 12'b000001000100;
		12'd728:BCD_Out <= 12'b000001000100;
		12'd729:BCD_Out <= 12'b000001000101;
		12'd730:BCD_Out <= 12'b000001000101;
		12'd731:BCD_Out <= 12'b000001000101;
		12'd732:BCD_Out <= 12'b000001000101;
		12'd733:BCD_Out <= 12'b000001000101;
		12'd734:BCD_Out <= 12'b000001000101;
		12'd735:BCD_Out <= 12'b000001000101;
		12'd736:BCD_Out <= 12'b000001000101;
		12'd737:BCD_Out <= 12'b000001000101;
		12'd738:BCD_Out <= 12'b000001000101;
		12'd739:BCD_Out <= 12'b000001000101;
		12'd740:BCD_Out <= 12'b000001000101;
		12'd741:BCD_Out <= 12'b000001000101;
		12'd742:BCD_Out <= 12'b000001000101;
		12'd743:BCD_Out <= 12'b000001000101;
		12'd744:BCD_Out <= 12'b000001000101;
		12'd745:BCD_Out <= 12'b000001000101;
		12'd746:BCD_Out <= 12'b000001000110;
		12'd747:BCD_Out <= 12'b000001000110;
		12'd748:BCD_Out <= 12'b000001000110;
		12'd749:BCD_Out <= 12'b000001000110;
		12'd750:BCD_Out <= 12'b000001000110;
		12'd751:BCD_Out <= 12'b000001000110;
		12'd752:BCD_Out <= 12'b000001000110;
		12'd753:BCD_Out <= 12'b000001000110;
		12'd754:BCD_Out <= 12'b000001000110;
		12'd755:BCD_Out <= 12'b000001000110;
		12'd756:BCD_Out <= 12'b000001000110;
		12'd757:BCD_Out <= 12'b000001000110;
		12'd758:BCD_Out <= 12'b000001000110;
		12'd759:BCD_Out <= 12'b000001000110;
		12'd760:BCD_Out <= 12'b000001000110;
		12'd761:BCD_Out <= 12'b000001000110;
		12'd762:BCD_Out <= 12'b000001000111;
		12'd763:BCD_Out <= 12'b000001000111;
		12'd764:BCD_Out <= 12'b000001000111;
		12'd765:BCD_Out <= 12'b000001000111;
		12'd766:BCD_Out <= 12'b000001000111;
		12'd767:BCD_Out <= 12'b000001000111;
		12'd768:BCD_Out <= 12'b000001000111;
		12'd769:BCD_Out <= 12'b000001000111;
		12'd770:BCD_Out <= 12'b000001000111;
		12'd771:BCD_Out <= 12'b000001000111;
		12'd772:BCD_Out <= 12'b000001000111;
		12'd773:BCD_Out <= 12'b000001000111;
		12'd774:BCD_Out <= 12'b000001000111;
		12'd775:BCD_Out <= 12'b000001000111;
		12'd776:BCD_Out <= 12'b000001000111;
		12'd777:BCD_Out <= 12'b000001000111;
		12'd778:BCD_Out <= 12'b000001000111;
		12'd779:BCD_Out <= 12'b000001001000;
		12'd780:BCD_Out <= 12'b000001001000;
		12'd781:BCD_Out <= 12'b000001001000;
		12'd782:BCD_Out <= 12'b000001001000;
		12'd783:BCD_Out <= 12'b000001001000;
		12'd784:BCD_Out <= 12'b000001001000;
		12'd785:BCD_Out <= 12'b000001001000;
		12'd786:BCD_Out <= 12'b000001001000;
		12'd787:BCD_Out <= 12'b000001001000;
		12'd788:BCD_Out <= 12'b000001001000;
		12'd789:BCD_Out <= 12'b000001001000;
		12'd790:BCD_Out <= 12'b000001001000;
		12'd791:BCD_Out <= 12'b000001001000;
		12'd792:BCD_Out <= 12'b000001001000;
		12'd793:BCD_Out <= 12'b000001001000;
		12'd794:BCD_Out <= 12'b000001001000;
		12'd795:BCD_Out <= 12'b000001001001;
		12'd796:BCD_Out <= 12'b000001001001;
		12'd797:BCD_Out <= 12'b000001001001;
		12'd798:BCD_Out <= 12'b000001001001;
		12'd799:BCD_Out <= 12'b000001001001;
		12'd800:BCD_Out <= 12'b000001001001;
		12'd801:BCD_Out <= 12'b000001001001;
		12'd802:BCD_Out <= 12'b000001001001;
		12'd803:BCD_Out <= 12'b000001001001;
		12'd804:BCD_Out <= 12'b000001001001;
		12'd805:BCD_Out <= 12'b000001001001;
		12'd806:BCD_Out <= 12'b000001001001;
		12'd807:BCD_Out <= 12'b000001001001;
		12'd808:BCD_Out <= 12'b000001001001;
		12'd809:BCD_Out <= 12'b000001001001;
		12'd810:BCD_Out <= 12'b000001001001;
		12'd811:BCD_Out <= 12'b000001010000;
		12'd812:BCD_Out <= 12'b000001010000;
		12'd813:BCD_Out <= 12'b000001010000;
		12'd814:BCD_Out <= 12'b000001010000;
		12'd815:BCD_Out <= 12'b000001010000;
		12'd816:BCD_Out <= 12'b000001010000;
		12'd817:BCD_Out <= 12'b000001010000;
		12'd818:BCD_Out <= 12'b000001010000;
		12'd819:BCD_Out <= 12'b000001010000;
		12'd820:BCD_Out <= 12'b000001010000;
		12'd821:BCD_Out <= 12'b000001010000;
		12'd822:BCD_Out <= 12'b000001010000;
		12'd823:BCD_Out <= 12'b000001010000;
		12'd824:BCD_Out <= 12'b000001010000;
		12'd825:BCD_Out <= 12'b000001010000;
		12'd826:BCD_Out <= 12'b000001010000;
		12'd827:BCD_Out <= 12'b000001010000;
		12'd828:BCD_Out <= 12'b000001010001;
		12'd829:BCD_Out <= 12'b000001010001;
		12'd830:BCD_Out <= 12'b000001010001;
		12'd831:BCD_Out <= 12'b000001010001;
		12'd832:BCD_Out <= 12'b000001010001;
		12'd833:BCD_Out <= 12'b000001010001;
		12'd834:BCD_Out <= 12'b000001010001;
		12'd835:BCD_Out <= 12'b000001010001;
		12'd836:BCD_Out <= 12'b000001010001;
		12'd837:BCD_Out <= 12'b000001010001;
		12'd838:BCD_Out <= 12'b000001010001;
		12'd839:BCD_Out <= 12'b000001010001;
		12'd840:BCD_Out <= 12'b000001010001;
		12'd841:BCD_Out <= 12'b000001010001;
		12'd842:BCD_Out <= 12'b000001010001;
		12'd843:BCD_Out <= 12'b000001010001;
		12'd844:BCD_Out <= 12'b000001010010;
		12'd845:BCD_Out <= 12'b000001010010;
		12'd846:BCD_Out <= 12'b000001010010;
		12'd847:BCD_Out <= 12'b000001010010;
		12'd848:BCD_Out <= 12'b000001010010;
		12'd849:BCD_Out <= 12'b000001010010;
		12'd850:BCD_Out <= 12'b000001010010;
		12'd851:BCD_Out <= 12'b000001010010;
		12'd852:BCD_Out <= 12'b000001010010;
		12'd853:BCD_Out <= 12'b000001010010;
		12'd854:BCD_Out <= 12'b000001010010;
		12'd855:BCD_Out <= 12'b000001010010;
		12'd856:BCD_Out <= 12'b000001010010;
		12'd857:BCD_Out <= 12'b000001010010;
		12'd858:BCD_Out <= 12'b000001010010;
		12'd859:BCD_Out <= 12'b000001010010;
		12'd860:BCD_Out <= 12'b000001010011;
		12'd861:BCD_Out <= 12'b000001010011;
		12'd862:BCD_Out <= 12'b000001010011;
		12'd863:BCD_Out <= 12'b000001010011;
		12'd864:BCD_Out <= 12'b000001010011;
		12'd865:BCD_Out <= 12'b000001010011;
		12'd866:BCD_Out <= 12'b000001010011;
		12'd867:BCD_Out <= 12'b000001010011;
		12'd868:BCD_Out <= 12'b000001010011;
		12'd869:BCD_Out <= 12'b000001010011;
		12'd870:BCD_Out <= 12'b000001010011;
		12'd871:BCD_Out <= 12'b000001010011;
		12'd872:BCD_Out <= 12'b000001010011;
		12'd873:BCD_Out <= 12'b000001010011;
		12'd874:BCD_Out <= 12'b000001010011;
		12'd875:BCD_Out <= 12'b000001010011;
		12'd876:BCD_Out <= 12'b000001010011;
		12'd877:BCD_Out <= 12'b000001010100;
		12'd878:BCD_Out <= 12'b000001010100;
		12'd879:BCD_Out <= 12'b000001010100;
		12'd880:BCD_Out <= 12'b000001010100;
		12'd881:BCD_Out <= 12'b000001010100;
		12'd882:BCD_Out <= 12'b000001010100;
		12'd883:BCD_Out <= 12'b000001010100;
		12'd884:BCD_Out <= 12'b000001010100;
		12'd885:BCD_Out <= 12'b000001010100;
		12'd886:BCD_Out <= 12'b000001010100;
		12'd887:BCD_Out <= 12'b000001010100;
		12'd888:BCD_Out <= 12'b000001010100;
		12'd889:BCD_Out <= 12'b000001010100;
		12'd890:BCD_Out <= 12'b000001010100;
		12'd891:BCD_Out <= 12'b000001010100;
		12'd892:BCD_Out <= 12'b000001010100;
		12'd893:BCD_Out <= 12'b000001010101;
		12'd894:BCD_Out <= 12'b000001010101;
		12'd895:BCD_Out <= 12'b000001010101;
		12'd896:BCD_Out <= 12'b000001010101;
		12'd897:BCD_Out <= 12'b000001010101;
		12'd898:BCD_Out <= 12'b000001010101;
		12'd899:BCD_Out <= 12'b000001010101;
		12'd900:BCD_Out <= 12'b000001010101;
		12'd901:BCD_Out <= 12'b000001010101;
		12'd902:BCD_Out <= 12'b000001010101;
		12'd903:BCD_Out <= 12'b000001010101;
		12'd904:BCD_Out <= 12'b000001010101;
		12'd905:BCD_Out <= 12'b000001010101;
		12'd906:BCD_Out <= 12'b000001010101;
		12'd907:BCD_Out <= 12'b000001010101;
		12'd908:BCD_Out <= 12'b000001010101;
		12'd909:BCD_Out <= 12'b000001010101;
		12'd910:BCD_Out <= 12'b000001010110;
		12'd911:BCD_Out <= 12'b000001010110;
		12'd912:BCD_Out <= 12'b000001010110;
		12'd913:BCD_Out <= 12'b000001010110;
		12'd914:BCD_Out <= 12'b000001010110;
		12'd915:BCD_Out <= 12'b000001010110;
		12'd916:BCD_Out <= 12'b000001010110;
		12'd917:BCD_Out <= 12'b000001010110;
		12'd918:BCD_Out <= 12'b000001010110;
		12'd919:BCD_Out <= 12'b000001010110;
		12'd920:BCD_Out <= 12'b000001010110;
		12'd921:BCD_Out <= 12'b000001010110;
		12'd922:BCD_Out <= 12'b000001010110;
		12'd923:BCD_Out <= 12'b000001010110;
		12'd924:BCD_Out <= 12'b000001010110;
		12'd925:BCD_Out <= 12'b000001010110;
		12'd926:BCD_Out <= 12'b000001010111;
		12'd927:BCD_Out <= 12'b000001010111;
		12'd928:BCD_Out <= 12'b000001010111;
		12'd929:BCD_Out <= 12'b000001010111;
		12'd930:BCD_Out <= 12'b000001010111;
		12'd931:BCD_Out <= 12'b000001010111;
		12'd932:BCD_Out <= 12'b000001010111;
		12'd933:BCD_Out <= 12'b000001010111;
		12'd934:BCD_Out <= 12'b000001010111;
		12'd935:BCD_Out <= 12'b000001010111;
		12'd936:BCD_Out <= 12'b000001010111;
		12'd937:BCD_Out <= 12'b000001010111;
		12'd938:BCD_Out <= 12'b000001010111;
		12'd939:BCD_Out <= 12'b000001010111;
		12'd940:BCD_Out <= 12'b000001010111;
		12'd941:BCD_Out <= 12'b000001010111;
		12'd942:BCD_Out <= 12'b000001011000;
		12'd943:BCD_Out <= 12'b000001011000;
		12'd944:BCD_Out <= 12'b000001011000;
		12'd945:BCD_Out <= 12'b000001011000;
		12'd946:BCD_Out <= 12'b000001011000;
		12'd947:BCD_Out <= 12'b000001011000;
		12'd948:BCD_Out <= 12'b000001011000;
		12'd949:BCD_Out <= 12'b000001011000;
		12'd950:BCD_Out <= 12'b000001011000;
		12'd951:BCD_Out <= 12'b000001011000;
		12'd952:BCD_Out <= 12'b000001011000;
		12'd953:BCD_Out <= 12'b000001011000;
		12'd954:BCD_Out <= 12'b000001011000;
		12'd955:BCD_Out <= 12'b000001011000;
		12'd956:BCD_Out <= 12'b000001011000;
		12'd957:BCD_Out <= 12'b000001011000;
		12'd958:BCD_Out <= 12'b000001011000;
		12'd959:BCD_Out <= 12'b000001011001;
		12'd960:BCD_Out <= 12'b000001011001;
		12'd961:BCD_Out <= 12'b000001011001;
		12'd962:BCD_Out <= 12'b000001011001;
		12'd963:BCD_Out <= 12'b000001011001;
		12'd964:BCD_Out <= 12'b000001011001;
		12'd965:BCD_Out <= 12'b000001011001;
		12'd966:BCD_Out <= 12'b000001011001;
		12'd967:BCD_Out <= 12'b000001011001;
		12'd968:BCD_Out <= 12'b000001011001;
		12'd969:BCD_Out <= 12'b000001011001;
		12'd970:BCD_Out <= 12'b000001011001;
		12'd971:BCD_Out <= 12'b000001011001;
		12'd972:BCD_Out <= 12'b000001011001;
		12'd973:BCD_Out <= 12'b000001011001;
		12'd974:BCD_Out <= 12'b000001011001;
		12'd975:BCD_Out <= 12'b000001100000;
		12'd976:BCD_Out <= 12'b000001100000;
		12'd977:BCD_Out <= 12'b000001100000;
		12'd978:BCD_Out <= 12'b000001100000;
		12'd979:BCD_Out <= 12'b000001100000;
		12'd980:BCD_Out <= 12'b000001100000;
		12'd981:BCD_Out <= 12'b000001100000;
		12'd982:BCD_Out <= 12'b000001100000;
		12'd983:BCD_Out <= 12'b000001100000;
		12'd984:BCD_Out <= 12'b000001100000;
		12'd985:BCD_Out <= 12'b000001100000;
		12'd986:BCD_Out <= 12'b000001100000;
		12'd987:BCD_Out <= 12'b000001100000;
		12'd988:BCD_Out <= 12'b000001100000;
		12'd989:BCD_Out <= 12'b000001100000;
		12'd990:BCD_Out <= 12'b000001100000;
		12'd991:BCD_Out <= 12'b000001100001;
		12'd992:BCD_Out <= 12'b000001100001;
		12'd993:BCD_Out <= 12'b000001100001;
		12'd994:BCD_Out <= 12'b000001100001;
		12'd995:BCD_Out <= 12'b000001100001;
		12'd996:BCD_Out <= 12'b000001100001;
		12'd997:BCD_Out <= 12'b000001100001;
		12'd998:BCD_Out <= 12'b000001100001;
		12'd999:BCD_Out <= 12'b000001100001;
		12'd1000:BCD_Out <= 12'b000001100001;
		12'd1001:BCD_Out <= 12'b000001100001;
		12'd1002:BCD_Out <= 12'b000001100001;
		12'd1003:BCD_Out <= 12'b000001100001;
		12'd1004:BCD_Out <= 12'b000001100001;
		12'd1005:BCD_Out <= 12'b000001100001;
		12'd1006:BCD_Out <= 12'b000001100001;
		12'd1007:BCD_Out <= 12'b000001100001;
		12'd1008:BCD_Out <= 12'b000001100010;
		12'd1009:BCD_Out <= 12'b000001100010;
		12'd1010:BCD_Out <= 12'b000001100010;
		12'd1011:BCD_Out <= 12'b000001100010;
		12'd1012:BCD_Out <= 12'b000001100010;
		12'd1013:BCD_Out <= 12'b000001100010;
		12'd1014:BCD_Out <= 12'b000001100010;
		12'd1015:BCD_Out <= 12'b000001100010;
		12'd1016:BCD_Out <= 12'b000001100010;
		12'd1017:BCD_Out <= 12'b000001100010;
		12'd1018:BCD_Out <= 12'b000001100010;
		12'd1019:BCD_Out <= 12'b000001100010;
		12'd1020:BCD_Out <= 12'b000001100010;
		12'd1021:BCD_Out <= 12'b000001100010;
		12'd1022:BCD_Out <= 12'b000001100010;
		12'd1023:BCD_Out <= 12'b000001100010;
		12'd1024:BCD_Out <= 12'b000001100011;
		12'd1025:BCD_Out <= 12'b000001100011;
		12'd1026:BCD_Out <= 12'b000001100011;
		12'd1027:BCD_Out <= 12'b000001100011;
		12'd1028:BCD_Out <= 12'b000001100011;
		12'd1029:BCD_Out <= 12'b000001100011;
		12'd1030:BCD_Out <= 12'b000001100011;
		12'd1031:BCD_Out <= 12'b000001100011;
		12'd1032:BCD_Out <= 12'b000001100011;
		12'd1033:BCD_Out <= 12'b000001100011;
		12'd1034:BCD_Out <= 12'b000001100011;
		12'd1035:BCD_Out <= 12'b000001100011;
		12'd1036:BCD_Out <= 12'b000001100011;
		12'd1037:BCD_Out <= 12'b000001100011;
		12'd1038:BCD_Out <= 12'b000001100011;
		12'd1039:BCD_Out <= 12'b000001100011;
		12'd1040:BCD_Out <= 12'b000001100011;
		12'd1041:BCD_Out <= 12'b000001100100;
		12'd1042:BCD_Out <= 12'b000001100100;
		12'd1043:BCD_Out <= 12'b000001100100;
		12'd1044:BCD_Out <= 12'b000001100100;
		12'd1045:BCD_Out <= 12'b000001100100;
		12'd1046:BCD_Out <= 12'b000001100100;
		12'd1047:BCD_Out <= 12'b000001100100;
		12'd1048:BCD_Out <= 12'b000001100100;
		12'd1049:BCD_Out <= 12'b000001100100;
		12'd1050:BCD_Out <= 12'b000001100100;
		12'd1051:BCD_Out <= 12'b000001100100;
		12'd1052:BCD_Out <= 12'b000001100100;
		12'd1053:BCD_Out <= 12'b000001100100;
		12'd1054:BCD_Out <= 12'b000001100100;
		12'd1055:BCD_Out <= 12'b000001100100;
		12'd1056:BCD_Out <= 12'b000001100100;
		12'd1057:BCD_Out <= 12'b000001100101;
		12'd1058:BCD_Out <= 12'b000001100101;
		12'd1059:BCD_Out <= 12'b000001100101;
		12'd1060:BCD_Out <= 12'b000001100101;
		12'd1061:BCD_Out <= 12'b000001100101;
		12'd1062:BCD_Out <= 12'b000001100101;
		12'd1063:BCD_Out <= 12'b000001100101;
		12'd1064:BCD_Out <= 12'b000001100101;
		12'd1065:BCD_Out <= 12'b000001100101;
		12'd1066:BCD_Out <= 12'b000001100101;
		12'd1067:BCD_Out <= 12'b000001100101;
		12'd1068:BCD_Out <= 12'b000001100101;
		12'd1069:BCD_Out <= 12'b000001100101;
		12'd1070:BCD_Out <= 12'b000001100101;
		12'd1071:BCD_Out <= 12'b000001100101;
		12'd1072:BCD_Out <= 12'b000001100101;
		12'd1073:BCD_Out <= 12'b000001100110;
		12'd1074:BCD_Out <= 12'b000001100110;
		12'd1075:BCD_Out <= 12'b000001100110;
		12'd1076:BCD_Out <= 12'b000001100110;
		12'd1077:BCD_Out <= 12'b000001100110;
		12'd1078:BCD_Out <= 12'b000001100110;
		12'd1079:BCD_Out <= 12'b000001100110;
		12'd1080:BCD_Out <= 12'b000001100110;
		12'd1081:BCD_Out <= 12'b000001100110;
		12'd1082:BCD_Out <= 12'b000001100110;
		12'd1083:BCD_Out <= 12'b000001100110;
		12'd1084:BCD_Out <= 12'b000001100110;
		12'd1085:BCD_Out <= 12'b000001100110;
		12'd1086:BCD_Out <= 12'b000001100110;
		12'd1087:BCD_Out <= 12'b000001100110;
		12'd1088:BCD_Out <= 12'b000001100110;
		12'd1089:BCD_Out <= 12'b000001100110;
		12'd1090:BCD_Out <= 12'b000001100111;
		12'd1091:BCD_Out <= 12'b000001100111;
		12'd1092:BCD_Out <= 12'b000001100111;
		12'd1093:BCD_Out <= 12'b000001100111;
		12'd1094:BCD_Out <= 12'b000001100111;
		12'd1095:BCD_Out <= 12'b000001100111;
		12'd1096:BCD_Out <= 12'b000001100111;
		12'd1097:BCD_Out <= 12'b000001100111;
		12'd1098:BCD_Out <= 12'b000001100111;
		12'd1099:BCD_Out <= 12'b000001100111;
		12'd1100:BCD_Out <= 12'b000001100111;
		12'd1101:BCD_Out <= 12'b000001100111;
		12'd1102:BCD_Out <= 12'b000001100111;
		12'd1103:BCD_Out <= 12'b000001100111;
		12'd1104:BCD_Out <= 12'b000001100111;
		12'd1105:BCD_Out <= 12'b000001100111;
		12'd1106:BCD_Out <= 12'b000001101000;
		12'd1107:BCD_Out <= 12'b000001101000;
		12'd1108:BCD_Out <= 12'b000001101000;
		12'd1109:BCD_Out <= 12'b000001101000;
		12'd1110:BCD_Out <= 12'b000001101000;
		12'd1111:BCD_Out <= 12'b000001101000;
		12'd1112:BCD_Out <= 12'b000001101000;
		12'd1113:BCD_Out <= 12'b000001101000;
		12'd1114:BCD_Out <= 12'b000001101000;
		12'd1115:BCD_Out <= 12'b000001101000;
		12'd1116:BCD_Out <= 12'b000001101000;
		12'd1117:BCD_Out <= 12'b000001101000;
		12'd1118:BCD_Out <= 12'b000001101000;
		12'd1119:BCD_Out <= 12'b000001101000;
		12'd1120:BCD_Out <= 12'b000001101000;
		12'd1121:BCD_Out <= 12'b000001101000;
		12'd1122:BCD_Out <= 12'b000001101000;
		12'd1123:BCD_Out <= 12'b000001101001;
		12'd1124:BCD_Out <= 12'b000001101001;
		12'd1125:BCD_Out <= 12'b000001101001;
		12'd1126:BCD_Out <= 12'b000001101001;
		12'd1127:BCD_Out <= 12'b000001101001;
		12'd1128:BCD_Out <= 12'b000001101001;
		12'd1129:BCD_Out <= 12'b000001101001;
		12'd1130:BCD_Out <= 12'b000001101001;
		12'd1131:BCD_Out <= 12'b000001101001;
		12'd1132:BCD_Out <= 12'b000001101001;
		12'd1133:BCD_Out <= 12'b000001101001;
		12'd1134:BCD_Out <= 12'b000001101001;
		12'd1135:BCD_Out <= 12'b000001101001;
		12'd1136:BCD_Out <= 12'b000001101001;
		12'd1137:BCD_Out <= 12'b000001101001;
		12'd1138:BCD_Out <= 12'b000001101001;
		12'd1139:BCD_Out <= 12'b000001110000;
		12'd1140:BCD_Out <= 12'b000001110000;
		12'd1141:BCD_Out <= 12'b000001110000;
		12'd1142:BCD_Out <= 12'b000001110000;
		12'd1143:BCD_Out <= 12'b000001110000;
		12'd1144:BCD_Out <= 12'b000001110000;
		12'd1145:BCD_Out <= 12'b000001110000;
		12'd1146:BCD_Out <= 12'b000001110000;
		12'd1147:BCD_Out <= 12'b000001110000;
		12'd1148:BCD_Out <= 12'b000001110000;
		12'd1149:BCD_Out <= 12'b000001110000;
		12'd1150:BCD_Out <= 12'b000001110000;
		12'd1151:BCD_Out <= 12'b000001110000;
		12'd1152:BCD_Out <= 12'b000001110000;
		12'd1153:BCD_Out <= 12'b000001110000;
		12'd1154:BCD_Out <= 12'b000001110000;
		12'd1155:BCD_Out <= 12'b000001110001;
		12'd1156:BCD_Out <= 12'b000001110001;
		12'd1157:BCD_Out <= 12'b000001110001;
		12'd1158:BCD_Out <= 12'b000001110001;
		12'd1159:BCD_Out <= 12'b000001110001;
		12'd1160:BCD_Out <= 12'b000001110001;
		12'd1161:BCD_Out <= 12'b000001110001;
		12'd1162:BCD_Out <= 12'b000001110001;
		12'd1163:BCD_Out <= 12'b000001110001;
		12'd1164:BCD_Out <= 12'b000001110001;
		12'd1165:BCD_Out <= 12'b000001110001;
		12'd1166:BCD_Out <= 12'b000001110001;
		12'd1167:BCD_Out <= 12'b000001110001;
		12'd1168:BCD_Out <= 12'b000001110001;
		12'd1169:BCD_Out <= 12'b000001110001;
		12'd1170:BCD_Out <= 12'b000001110001;
		12'd1171:BCD_Out <= 12'b000001110001;
		12'd1172:BCD_Out <= 12'b000001110010;
		12'd1173:BCD_Out <= 12'b000001110010;
		12'd1174:BCD_Out <= 12'b000001110010;
		12'd1175:BCD_Out <= 12'b000001110010;
		12'd1176:BCD_Out <= 12'b000001110010;
		12'd1177:BCD_Out <= 12'b000001110010;
		12'd1178:BCD_Out <= 12'b000001110010;
		12'd1179:BCD_Out <= 12'b000001110010;
		12'd1180:BCD_Out <= 12'b000001110010;
		12'd1181:BCD_Out <= 12'b000001110010;
		12'd1182:BCD_Out <= 12'b000001110010;
		12'd1183:BCD_Out <= 12'b000001110010;
		12'd1184:BCD_Out <= 12'b000001110010;
		12'd1185:BCD_Out <= 12'b000001110010;
		12'd1186:BCD_Out <= 12'b000001110010;
		12'd1187:BCD_Out <= 12'b000001110010;
		12'd1188:BCD_Out <= 12'b000001110011;
		12'd1189:BCD_Out <= 12'b000001110011;
		12'd1190:BCD_Out <= 12'b000001110011;
		12'd1191:BCD_Out <= 12'b000001110011;
		12'd1192:BCD_Out <= 12'b000001110011;
		12'd1193:BCD_Out <= 12'b000001110011;
		12'd1194:BCD_Out <= 12'b000001110011;
		12'd1195:BCD_Out <= 12'b000001110011;
		12'd1196:BCD_Out <= 12'b000001110011;
		12'd1197:BCD_Out <= 12'b000001110011;
		12'd1198:BCD_Out <= 12'b000001110011;
		12'd1199:BCD_Out <= 12'b000001110011;
		12'd1200:BCD_Out <= 12'b000001110011;
		12'd1201:BCD_Out <= 12'b000001110011;
		12'd1202:BCD_Out <= 12'b000001110011;
		12'd1203:BCD_Out <= 12'b000001110011;
		12'd1204:BCD_Out <= 12'b000001110100;
		12'd1205:BCD_Out <= 12'b000001110100;
		12'd1206:BCD_Out <= 12'b000001110100;
		12'd1207:BCD_Out <= 12'b000001110100;
		12'd1208:BCD_Out <= 12'b000001110100;
		12'd1209:BCD_Out <= 12'b000001110100;
		12'd1210:BCD_Out <= 12'b000001110100;
		12'd1211:BCD_Out <= 12'b000001110100;
		12'd1212:BCD_Out <= 12'b000001110100;
		12'd1213:BCD_Out <= 12'b000001110100;
		12'd1214:BCD_Out <= 12'b000001110100;
		12'd1215:BCD_Out <= 12'b000001110100;
		12'd1216:BCD_Out <= 12'b000001110100;
		12'd1217:BCD_Out <= 12'b000001110100;
		12'd1218:BCD_Out <= 12'b000001110100;
		12'd1219:BCD_Out <= 12'b000001110100;
		12'd1220:BCD_Out <= 12'b000001110100;
		12'd1221:BCD_Out <= 12'b000001110101;
		12'd1222:BCD_Out <= 12'b000001110101;
		12'd1223:BCD_Out <= 12'b000001110101;
		12'd1224:BCD_Out <= 12'b000001110101;
		12'd1225:BCD_Out <= 12'b000001110101;
		12'd1226:BCD_Out <= 12'b000001110101;
		12'd1227:BCD_Out <= 12'b000001110101;
		12'd1228:BCD_Out <= 12'b000001110101;
		12'd1229:BCD_Out <= 12'b000001110101;
		12'd1230:BCD_Out <= 12'b000001110101;
		12'd1231:BCD_Out <= 12'b000001110101;
		12'd1232:BCD_Out <= 12'b000001110101;
		12'd1233:BCD_Out <= 12'b000001110101;
		12'd1234:BCD_Out <= 12'b000001110101;
		12'd1235:BCD_Out <= 12'b000001110101;
		12'd1236:BCD_Out <= 12'b000001110101;
		12'd1237:BCD_Out <= 12'b000001110110;
		12'd1238:BCD_Out <= 12'b000001110110;
		12'd1239:BCD_Out <= 12'b000001110110;
		12'd1240:BCD_Out <= 12'b000001110110;
		12'd1241:BCD_Out <= 12'b000001110110;
		12'd1242:BCD_Out <= 12'b000001110110;
		12'd1243:BCD_Out <= 12'b000001110110;
		12'd1244:BCD_Out <= 12'b000001110110;
		12'd1245:BCD_Out <= 12'b000001110110;
		12'd1246:BCD_Out <= 12'b000001110110;
		12'd1247:BCD_Out <= 12'b000001110110;
		12'd1248:BCD_Out <= 12'b000001110110;
		12'd1249:BCD_Out <= 12'b000001110110;
		12'd1250:BCD_Out <= 12'b000001110110;
		12'd1251:BCD_Out <= 12'b000001110110;
		12'd1252:BCD_Out <= 12'b000001110110;
		12'd1253:BCD_Out <= 12'b000001110110;
		12'd1254:BCD_Out <= 12'b000001110111;
		12'd1255:BCD_Out <= 12'b000001110111;
		12'd1256:BCD_Out <= 12'b000001110111;
		12'd1257:BCD_Out <= 12'b000001110111;
		12'd1258:BCD_Out <= 12'b000001110111;
		12'd1259:BCD_Out <= 12'b000001110111;
		12'd1260:BCD_Out <= 12'b000001110111;
		12'd1261:BCD_Out <= 12'b000001110111;
		12'd1262:BCD_Out <= 12'b000001110111;
		12'd1263:BCD_Out <= 12'b000001110111;
		12'd1264:BCD_Out <= 12'b000001110111;
		12'd1265:BCD_Out <= 12'b000001110111;
		12'd1266:BCD_Out <= 12'b000001110111;
		12'd1267:BCD_Out <= 12'b000001110111;
		12'd1268:BCD_Out <= 12'b000001110111;
		12'd1269:BCD_Out <= 12'b000001110111;
		12'd1270:BCD_Out <= 12'b000001111000;
		12'd1271:BCD_Out <= 12'b000001111000;
		12'd1272:BCD_Out <= 12'b000001111000;
		12'd1273:BCD_Out <= 12'b000001111000;
		12'd1274:BCD_Out <= 12'b000001111000;
		12'd1275:BCD_Out <= 12'b000001111000;
		12'd1276:BCD_Out <= 12'b000001111000;
		12'd1277:BCD_Out <= 12'b000001111000;
		12'd1278:BCD_Out <= 12'b000001111000;
		12'd1279:BCD_Out <= 12'b000001111000;
		12'd1280:BCD_Out <= 12'b000001111000;
		12'd1281:BCD_Out <= 12'b000001111000;
		12'd1282:BCD_Out <= 12'b000001111000;
		12'd1283:BCD_Out <= 12'b000001111000;
		12'd1284:BCD_Out <= 12'b000001111000;
		12'd1285:BCD_Out <= 12'b000001111000;
		12'd1286:BCD_Out <= 12'b000001111001;
		12'd1287:BCD_Out <= 12'b000001111001;
		12'd1288:BCD_Out <= 12'b000001111001;
		12'd1289:BCD_Out <= 12'b000001111001;
		12'd1290:BCD_Out <= 12'b000001111001;
		12'd1291:BCD_Out <= 12'b000001111001;
		12'd1292:BCD_Out <= 12'b000001111001;
		12'd1293:BCD_Out <= 12'b000001111001;
		12'd1294:BCD_Out <= 12'b000001111001;
		12'd1295:BCD_Out <= 12'b000001111001;
		12'd1296:BCD_Out <= 12'b000001111001;
		12'd1297:BCD_Out <= 12'b000001111001;
		12'd1298:BCD_Out <= 12'b000001111001;
		12'd1299:BCD_Out <= 12'b000001111001;
		12'd1300:BCD_Out <= 12'b000001111001;
		12'd1301:BCD_Out <= 12'b000001111001;
		12'd1302:BCD_Out <= 12'b000001111001;
		12'd1303:BCD_Out <= 12'b000010000000;
		12'd1304:BCD_Out <= 12'b000010000000;
		12'd1305:BCD_Out <= 12'b000010000000;
		12'd1306:BCD_Out <= 12'b000010000000;
		12'd1307:BCD_Out <= 12'b000010000000;
		12'd1308:BCD_Out <= 12'b000010000000;
		12'd1309:BCD_Out <= 12'b000010000000;
		12'd1310:BCD_Out <= 12'b000010000000;
		12'd1311:BCD_Out <= 12'b000010000000;
		12'd1312:BCD_Out <= 12'b000010000000;
		12'd1313:BCD_Out <= 12'b000010000000;
		12'd1314:BCD_Out <= 12'b000010000000;
		12'd1315:BCD_Out <= 12'b000010000000;
		12'd1316:BCD_Out <= 12'b000010000000;
		12'd1317:BCD_Out <= 12'b000010000000;
		12'd1318:BCD_Out <= 12'b000010000000;
		12'd1319:BCD_Out <= 12'b000010000001;
		12'd1320:BCD_Out <= 12'b000010000001;
		12'd1321:BCD_Out <= 12'b000010000001;
		12'd1322:BCD_Out <= 12'b000010000001;
		12'd1323:BCD_Out <= 12'b000010000001;
		12'd1324:BCD_Out <= 12'b000010000001;
		12'd1325:BCD_Out <= 12'b000010000001;
		12'd1326:BCD_Out <= 12'b000010000001;
		12'd1327:BCD_Out <= 12'b000010000001;
		12'd1328:BCD_Out <= 12'b000010000001;
		12'd1329:BCD_Out <= 12'b000010000001;
		12'd1330:BCD_Out <= 12'b000010000001;
		12'd1331:BCD_Out <= 12'b000010000001;
		12'd1332:BCD_Out <= 12'b000010000001;
		12'd1333:BCD_Out <= 12'b000010000001;
		12'd1334:BCD_Out <= 12'b000010000001;
		12'd1335:BCD_Out <= 12'b000010000010;
		12'd1336:BCD_Out <= 12'b000010000010;
		12'd1337:BCD_Out <= 12'b000010000010;
		12'd1338:BCD_Out <= 12'b000010000010;
		12'd1339:BCD_Out <= 12'b000010000010;
		12'd1340:BCD_Out <= 12'b000010000010;
		12'd1341:BCD_Out <= 12'b000010000010;
		12'd1342:BCD_Out <= 12'b000010000010;
		12'd1343:BCD_Out <= 12'b000010000010;
		12'd1344:BCD_Out <= 12'b000010000010;
		12'd1345:BCD_Out <= 12'b000010000010;
		12'd1346:BCD_Out <= 12'b000010000010;
		12'd1347:BCD_Out <= 12'b000010000010;
		12'd1348:BCD_Out <= 12'b000010000010;
		12'd1349:BCD_Out <= 12'b000010000010;
		12'd1350:BCD_Out <= 12'b000010000010;
		12'd1351:BCD_Out <= 12'b000010000010;
		12'd1352:BCD_Out <= 12'b000010000011;
		12'd1353:BCD_Out <= 12'b000010000011;
		12'd1354:BCD_Out <= 12'b000010000011;
		12'd1355:BCD_Out <= 12'b000010000011;
		12'd1356:BCD_Out <= 12'b000010000011;
		12'd1357:BCD_Out <= 12'b000010000011;
		12'd1358:BCD_Out <= 12'b000010000011;
		12'd1359:BCD_Out <= 12'b000010000011;
		12'd1360:BCD_Out <= 12'b000010000011;
		12'd1361:BCD_Out <= 12'b000010000011;
		12'd1362:BCD_Out <= 12'b000010000011;
		12'd1363:BCD_Out <= 12'b000010000011;
		12'd1364:BCD_Out <= 12'b000010000011;
		12'd1365:BCD_Out <= 12'b000010000011;
		12'd1366:BCD_Out <= 12'b000010000011;
		12'd1367:BCD_Out <= 12'b000010000011;
		12'd1368:BCD_Out <= 12'b000010000100;
		12'd1369:BCD_Out <= 12'b000010000100;
		12'd1370:BCD_Out <= 12'b000010000100;
		12'd1371:BCD_Out <= 12'b000010000100;
		12'd1372:BCD_Out <= 12'b000010000100;
		12'd1373:BCD_Out <= 12'b000010000100;
		12'd1374:BCD_Out <= 12'b000010000100;
		12'd1375:BCD_Out <= 12'b000010000100;
		12'd1376:BCD_Out <= 12'b000010000100;
		12'd1377:BCD_Out <= 12'b000010000100;
		12'd1378:BCD_Out <= 12'b000010000100;
		12'd1379:BCD_Out <= 12'b000010000100;
		12'd1380:BCD_Out <= 12'b000010000100;
		12'd1381:BCD_Out <= 12'b000010000100;
		12'd1382:BCD_Out <= 12'b000010000100;
		12'd1383:BCD_Out <= 12'b000010000100;
		12'd1384:BCD_Out <= 12'b000010000100;
		12'd1385:BCD_Out <= 12'b000010000101;
		12'd1386:BCD_Out <= 12'b000010000101;
		12'd1387:BCD_Out <= 12'b000010000101;
		12'd1388:BCD_Out <= 12'b000010000101;
		12'd1389:BCD_Out <= 12'b000010000101;
		12'd1390:BCD_Out <= 12'b000010000101;
		12'd1391:BCD_Out <= 12'b000010000101;
		12'd1392:BCD_Out <= 12'b000010000101;
		12'd1393:BCD_Out <= 12'b000010000101;
		12'd1394:BCD_Out <= 12'b000010000101;
		12'd1395:BCD_Out <= 12'b000010000101;
		12'd1396:BCD_Out <= 12'b000010000101;
		12'd1397:BCD_Out <= 12'b000010000101;
		12'd1398:BCD_Out <= 12'b000010000101;
		12'd1399:BCD_Out <= 12'b000010000101;
		12'd1400:BCD_Out <= 12'b000010000101;
		12'd1401:BCD_Out <= 12'b000010000110;
		12'd1402:BCD_Out <= 12'b000010000110;
		12'd1403:BCD_Out <= 12'b000010000110;
		12'd1404:BCD_Out <= 12'b000010000110;
		12'd1405:BCD_Out <= 12'b000010000110;
		12'd1406:BCD_Out <= 12'b000010000110;
		12'd1407:BCD_Out <= 12'b000010000110;
		12'd1408:BCD_Out <= 12'b000010000110;
		12'd1409:BCD_Out <= 12'b000010000110;
		12'd1410:BCD_Out <= 12'b000010000110;
		12'd1411:BCD_Out <= 12'b000010000110;
		12'd1412:BCD_Out <= 12'b000010000110;
		12'd1413:BCD_Out <= 12'b000010000110;
		12'd1414:BCD_Out <= 12'b000010000110;
		12'd1415:BCD_Out <= 12'b000010000110;
		12'd1416:BCD_Out <= 12'b000010000110;
		12'd1417:BCD_Out <= 12'b000010000111;
		12'd1418:BCD_Out <= 12'b000010000111;
		12'd1419:BCD_Out <= 12'b000010000111;
		12'd1420:BCD_Out <= 12'b000010000111;
		12'd1421:BCD_Out <= 12'b000010000111;
		12'd1422:BCD_Out <= 12'b000010000111;
		12'd1423:BCD_Out <= 12'b000010000111;
		12'd1424:BCD_Out <= 12'b000010000111;
		12'd1425:BCD_Out <= 12'b000010000111;
		12'd1426:BCD_Out <= 12'b000010000111;
		12'd1427:BCD_Out <= 12'b000010000111;
		12'd1428:BCD_Out <= 12'b000010000111;
		12'd1429:BCD_Out <= 12'b000010000111;
		12'd1430:BCD_Out <= 12'b000010000111;
		12'd1431:BCD_Out <= 12'b000010000111;
		12'd1432:BCD_Out <= 12'b000010000111;
		12'd1433:BCD_Out <= 12'b000010000111;
		12'd1434:BCD_Out <= 12'b000010001000;
		12'd1435:BCD_Out <= 12'b000010001000;
		12'd1436:BCD_Out <= 12'b000010001000;
		12'd1437:BCD_Out <= 12'b000010001000;
		12'd1438:BCD_Out <= 12'b000010001000;
		12'd1439:BCD_Out <= 12'b000010001000;
		12'd1440:BCD_Out <= 12'b000010001000;
		12'd1441:BCD_Out <= 12'b000010001000;
		12'd1442:BCD_Out <= 12'b000010001000;
		12'd1443:BCD_Out <= 12'b000010001000;
		12'd1444:BCD_Out <= 12'b000010001000;
		12'd1445:BCD_Out <= 12'b000010001000;
		12'd1446:BCD_Out <= 12'b000010001000;
		12'd1447:BCD_Out <= 12'b000010001000;
		12'd1448:BCD_Out <= 12'b000010001000;
		12'd1449:BCD_Out <= 12'b000010001000;
		12'd1450:BCD_Out <= 12'b000010001001;
		12'd1451:BCD_Out <= 12'b000010001001;
		12'd1452:BCD_Out <= 12'b000010001001;
		12'd1453:BCD_Out <= 12'b000010001001;
		12'd1454:BCD_Out <= 12'b000010001001;
		12'd1455:BCD_Out <= 12'b000010001001;
		12'd1456:BCD_Out <= 12'b000010001001;
		12'd1457:BCD_Out <= 12'b000010001001;
		12'd1458:BCD_Out <= 12'b000010001001;
		12'd1459:BCD_Out <= 12'b000010001001;
		12'd1460:BCD_Out <= 12'b000010001001;
		12'd1461:BCD_Out <= 12'b000010001001;
		12'd1462:BCD_Out <= 12'b000010001001;
		12'd1463:BCD_Out <= 12'b000010001001;
		12'd1464:BCD_Out <= 12'b000010001001;
		12'd1465:BCD_Out <= 12'b000010001001;
		12'd1466:BCD_Out <= 12'b000010001001;
		12'd1467:BCD_Out <= 12'b000010010000;
		12'd1468:BCD_Out <= 12'b000010010000;
		12'd1469:BCD_Out <= 12'b000010010000;
		12'd1470:BCD_Out <= 12'b000010010000;
		12'd1471:BCD_Out <= 12'b000010010000;
		12'd1472:BCD_Out <= 12'b000010010000;
		12'd1473:BCD_Out <= 12'b000010010000;
		12'd1474:BCD_Out <= 12'b000010010000;
		12'd1475:BCD_Out <= 12'b000010010000;
		12'd1476:BCD_Out <= 12'b000010010000;
		12'd1477:BCD_Out <= 12'b000010010000;
		12'd1478:BCD_Out <= 12'b000010010000;
		12'd1479:BCD_Out <= 12'b000010010000;
		12'd1480:BCD_Out <= 12'b000010010000;
		12'd1481:BCD_Out <= 12'b000010010000;
		12'd1482:BCD_Out <= 12'b000010010000;
		12'd1483:BCD_Out <= 12'b000010010001;
		12'd1484:BCD_Out <= 12'b000010010001;
		12'd1485:BCD_Out <= 12'b000010010001;
		12'd1486:BCD_Out <= 12'b000010010001;
		12'd1487:BCD_Out <= 12'b000010010001;
		12'd1488:BCD_Out <= 12'b000010010001;
		12'd1489:BCD_Out <= 12'b000010010001;
		12'd1490:BCD_Out <= 12'b000010010001;
		12'd1491:BCD_Out <= 12'b000010010001;
		12'd1492:BCD_Out <= 12'b000010010001;
		12'd1493:BCD_Out <= 12'b000010010001;
		12'd1494:BCD_Out <= 12'b000010010001;
		12'd1495:BCD_Out <= 12'b000010010001;
		12'd1496:BCD_Out <= 12'b000010010001;
		12'd1497:BCD_Out <= 12'b000010010001;
		12'd1498:BCD_Out <= 12'b000010010001;
		12'd1499:BCD_Out <= 12'b000010010010;
		12'd1500:BCD_Out <= 12'b000010010010;
		12'd1501:BCD_Out <= 12'b000010010010;
		12'd1502:BCD_Out <= 12'b000010010010;
		12'd1503:BCD_Out <= 12'b000010010010;
		12'd1504:BCD_Out <= 12'b000010010010;
		12'd1505:BCD_Out <= 12'b000010010010;
		12'd1506:BCD_Out <= 12'b000010010010;
		12'd1507:BCD_Out <= 12'b000010010010;
		12'd1508:BCD_Out <= 12'b000010010010;
		12'd1509:BCD_Out <= 12'b000010010010;
		12'd1510:BCD_Out <= 12'b000010010010;
		12'd1511:BCD_Out <= 12'b000010010010;
		12'd1512:BCD_Out <= 12'b000010010010;
		12'd1513:BCD_Out <= 12'b000010010010;
		12'd1514:BCD_Out <= 12'b000010010010;
		12'd1515:BCD_Out <= 12'b000010010010;
		12'd1516:BCD_Out <= 12'b000010010011;
		12'd1517:BCD_Out <= 12'b000010010011;
		12'd1518:BCD_Out <= 12'b000010010011;
		12'd1519:BCD_Out <= 12'b000010010011;
		12'd1520:BCD_Out <= 12'b000010010011;
		12'd1521:BCD_Out <= 12'b000010010011;
		12'd1522:BCD_Out <= 12'b000010010011;
		12'd1523:BCD_Out <= 12'b000010010011;
		12'd1524:BCD_Out <= 12'b000010010011;
		12'd1525:BCD_Out <= 12'b000010010011;
		12'd1526:BCD_Out <= 12'b000010010011;
		12'd1527:BCD_Out <= 12'b000010010011;
		12'd1528:BCD_Out <= 12'b000010010011;
		12'd1529:BCD_Out <= 12'b000010010011;
		12'd1530:BCD_Out <= 12'b000010010011;
		12'd1531:BCD_Out <= 12'b000010010011;
		12'd1532:BCD_Out <= 12'b000010010100;
		12'd1533:BCD_Out <= 12'b000010010100;
		12'd1534:BCD_Out <= 12'b000010010100;
		12'd1535:BCD_Out <= 12'b000010010100;
		12'd1536:BCD_Out <= 12'b000010010100;
		12'd1537:BCD_Out <= 12'b000010010100;
		12'd1538:BCD_Out <= 12'b000010010100;
		12'd1539:BCD_Out <= 12'b000010010100;
		12'd1540:BCD_Out <= 12'b000010010100;
		12'd1541:BCD_Out <= 12'b000010010100;
		12'd1542:BCD_Out <= 12'b000010010100;
		12'd1543:BCD_Out <= 12'b000010010100;
		12'd1544:BCD_Out <= 12'b000010010100;
		12'd1545:BCD_Out <= 12'b000010010100;
		12'd1546:BCD_Out <= 12'b000010010100;
		12'd1547:BCD_Out <= 12'b000010010100;
		12'd1548:BCD_Out <= 12'b000010010101;
		12'd1549:BCD_Out <= 12'b000010010101;
		12'd1550:BCD_Out <= 12'b000010010101;
		12'd1551:BCD_Out <= 12'b000010010101;
		12'd1552:BCD_Out <= 12'b000010010101;
		12'd1553:BCD_Out <= 12'b000010010101;
		12'd1554:BCD_Out <= 12'b000010010101;
		12'd1555:BCD_Out <= 12'b000010010101;
		12'd1556:BCD_Out <= 12'b000010010101;
		12'd1557:BCD_Out <= 12'b000010010101;
		12'd1558:BCD_Out <= 12'b000010010101;
		12'd1559:BCD_Out <= 12'b000010010101;
		12'd1560:BCD_Out <= 12'b000010010101;
		12'd1561:BCD_Out <= 12'b000010010101;
		12'd1562:BCD_Out <= 12'b000010010101;
		12'd1563:BCD_Out <= 12'b000010010101;
		12'd1564:BCD_Out <= 12'b000010010101;
		12'd1565:BCD_Out <= 12'b000010010110;
		12'd1566:BCD_Out <= 12'b000010010110;
		12'd1567:BCD_Out <= 12'b000010010110;
		12'd1568:BCD_Out <= 12'b000010010110;
		12'd1569:BCD_Out <= 12'b000010010110;
		12'd1570:BCD_Out <= 12'b000010010110;
		12'd1571:BCD_Out <= 12'b000010010110;
		12'd1572:BCD_Out <= 12'b000010010110;
		12'd1573:BCD_Out <= 12'b000010010110;
		12'd1574:BCD_Out <= 12'b000010010110;
		12'd1575:BCD_Out <= 12'b000010010110;
		12'd1576:BCD_Out <= 12'b000010010110;
		12'd1577:BCD_Out <= 12'b000010010110;
		12'd1578:BCD_Out <= 12'b000010010110;
		12'd1579:BCD_Out <= 12'b000010010110;
		12'd1580:BCD_Out <= 12'b000010010110;
		12'd1581:BCD_Out <= 12'b000010010111;
		12'd1582:BCD_Out <= 12'b000010010111;
		12'd1583:BCD_Out <= 12'b000010010111;
		12'd1584:BCD_Out <= 12'b000010010111;
		12'd1585:BCD_Out <= 12'b000010010111;
		12'd1586:BCD_Out <= 12'b000010010111;
		12'd1587:BCD_Out <= 12'b000010010111;
		12'd1588:BCD_Out <= 12'b000010010111;
		12'd1589:BCD_Out <= 12'b000010010111;
		12'd1590:BCD_Out <= 12'b000010010111;
		12'd1591:BCD_Out <= 12'b000010010111;
		12'd1592:BCD_Out <= 12'b000010010111;
		12'd1593:BCD_Out <= 12'b000010010111;
		12'd1594:BCD_Out <= 12'b000010010111;
		12'd1595:BCD_Out <= 12'b000010010111;
		12'd1596:BCD_Out <= 12'b000010010111;
		12'd1597:BCD_Out <= 12'b000010010111;
		12'd1598:BCD_Out <= 12'b000010011000;
		12'd1599:BCD_Out <= 12'b000010011000;
		12'd1600:BCD_Out <= 12'b000010011000;
		12'd1601:BCD_Out <= 12'b000010011000;
		12'd1602:BCD_Out <= 12'b000010011000;
		12'd1603:BCD_Out <= 12'b000010011000;
		12'd1604:BCD_Out <= 12'b000010011000;
		12'd1605:BCD_Out <= 12'b000010011000;
		12'd1606:BCD_Out <= 12'b000010011000;
		12'd1607:BCD_Out <= 12'b000010011000;
		12'd1608:BCD_Out <= 12'b000010011000;
		12'd1609:BCD_Out <= 12'b000010011000;
		12'd1610:BCD_Out <= 12'b000010011000;
		12'd1611:BCD_Out <= 12'b000010011000;
		12'd1612:BCD_Out <= 12'b000010011000;
		12'd1613:BCD_Out <= 12'b000010011000;
		12'd1614:BCD_Out <= 12'b000010011001;
		12'd1615:BCD_Out <= 12'b000010011001;
		12'd1616:BCD_Out <= 12'b000010011001;
		12'd1617:BCD_Out <= 12'b000010011001;
		12'd1618:BCD_Out <= 12'b000010011001;
		12'd1619:BCD_Out <= 12'b000010011001;
		12'd1620:BCD_Out <= 12'b000010011001;
		12'd1621:BCD_Out <= 12'b000010011001;
		12'd1622:BCD_Out <= 12'b000010011001;
		12'd1623:BCD_Out <= 12'b000010011001;
		12'd1624:BCD_Out <= 12'b000010011001;
		12'd1625:BCD_Out <= 12'b000010011001;
		12'd1626:BCD_Out <= 12'b000010011001;
		12'd1627:BCD_Out <= 12'b000010011001;
		12'd1628:BCD_Out <= 12'b000010011001;
		12'd1629:BCD_Out <= 12'b000010011001;
		12'd1630:BCD_Out <= 12'b000100000000;
		12'd1631:BCD_Out <= 12'b000100000000;
		12'd1632:BCD_Out <= 12'b000100000000;
		12'd1633:BCD_Out <= 12'b000100000000;
		12'd1634:BCD_Out <= 12'b000100000000;
		12'd1635:BCD_Out <= 12'b000100000000;
		12'd1636:BCD_Out <= 12'b000100000000;
		12'd1637:BCD_Out <= 12'b000100000000;
		12'd1638:BCD_Out <= 12'b000100000000;
		12'd1639:BCD_Out <= 12'b000100000000;
		12'd1640:BCD_Out <= 12'b000100000000;
		12'd1641:BCD_Out <= 12'b000100000000;
		12'd1642:BCD_Out <= 12'b000100000000;
		12'd1643:BCD_Out <= 12'b000100000000;
		12'd1644:BCD_Out <= 12'b000100000000;
		12'd1645:BCD_Out <= 12'b000100000000;
		12'd1646:BCD_Out <= 12'b000100000000;
		12'd1647:BCD_Out <= 12'b000100000001;
		12'd1648:BCD_Out <= 12'b000100000001;
		12'd1649:BCD_Out <= 12'b000100000001;
		12'd1650:BCD_Out <= 12'b000100000001;
		12'd1651:BCD_Out <= 12'b000100000001;
		12'd1652:BCD_Out <= 12'b000100000001;
		12'd1653:BCD_Out <= 12'b000100000001;
		12'd1654:BCD_Out <= 12'b000100000001;
		12'd1655:BCD_Out <= 12'b000100000001;
		12'd1656:BCD_Out <= 12'b000100000001;
		12'd1657:BCD_Out <= 12'b000100000001;
		12'd1658:BCD_Out <= 12'b000100000001;
		12'd1659:BCD_Out <= 12'b000100000001;
		12'd1660:BCD_Out <= 12'b000100000001;
		12'd1661:BCD_Out <= 12'b000100000001;
		12'd1662:BCD_Out <= 12'b000100000001;
		12'd1663:BCD_Out <= 12'b000100000010;
		12'd1664:BCD_Out <= 12'b000100000010;
		12'd1665:BCD_Out <= 12'b000100000010;
		12'd1666:BCD_Out <= 12'b000100000010;
		12'd1667:BCD_Out <= 12'b000100000010;
		12'd1668:BCD_Out <= 12'b000100000010;
		12'd1669:BCD_Out <= 12'b000100000010;
		12'd1670:BCD_Out <= 12'b000100000010;
		12'd1671:BCD_Out <= 12'b000100000010;
		12'd1672:BCD_Out <= 12'b000100000010;
		12'd1673:BCD_Out <= 12'b000100000010;
		12'd1674:BCD_Out <= 12'b000100000010;
		12'd1675:BCD_Out <= 12'b000100000010;
		12'd1676:BCD_Out <= 12'b000100000010;
		12'd1677:BCD_Out <= 12'b000100000010;
		12'd1678:BCD_Out <= 12'b000100000010;
		12'd1679:BCD_Out <= 12'b000100000011;
		12'd1680:BCD_Out <= 12'b000100000011;
		12'd1681:BCD_Out <= 12'b000100000011;
		12'd1682:BCD_Out <= 12'b000100000011;
		12'd1683:BCD_Out <= 12'b000100000011;
		12'd1684:BCD_Out <= 12'b000100000011;
		12'd1685:BCD_Out <= 12'b000100000011;
		12'd1686:BCD_Out <= 12'b000100000011;
		12'd1687:BCD_Out <= 12'b000100000011;
		12'd1688:BCD_Out <= 12'b000100000011;
		12'd1689:BCD_Out <= 12'b000100000011;
		12'd1690:BCD_Out <= 12'b000100000011;
		12'd1691:BCD_Out <= 12'b000100000011;
		12'd1692:BCD_Out <= 12'b000100000011;
		12'd1693:BCD_Out <= 12'b000100000011;
		12'd1694:BCD_Out <= 12'b000100000011;
		12'd1695:BCD_Out <= 12'b000100000011;
		12'd1696:BCD_Out <= 12'b000100000100;
		12'd1697:BCD_Out <= 12'b000100000100;
		12'd1698:BCD_Out <= 12'b000100000100;
		12'd1699:BCD_Out <= 12'b000100000100;
		12'd1700:BCD_Out <= 12'b000100000100;
		12'd1701:BCD_Out <= 12'b000100000100;
		12'd1702:BCD_Out <= 12'b000100000100;
		12'd1703:BCD_Out <= 12'b000100000100;
		12'd1704:BCD_Out <= 12'b000100000100;
		12'd1705:BCD_Out <= 12'b000100000100;
		12'd1706:BCD_Out <= 12'b000100000100;
		12'd1707:BCD_Out <= 12'b000100000100;
		12'd1708:BCD_Out <= 12'b000100000100;
		12'd1709:BCD_Out <= 12'b000100000100;
		12'd1710:BCD_Out <= 12'b000100000100;
		12'd1711:BCD_Out <= 12'b000100000100;
		12'd1712:BCD_Out <= 12'b000100000101;
		12'd1713:BCD_Out <= 12'b000100000101;
		12'd1714:BCD_Out <= 12'b000100000101;
		12'd1715:BCD_Out <= 12'b000100000101;
		12'd1716:BCD_Out <= 12'b000100000101;
		12'd1717:BCD_Out <= 12'b000100000101;
		12'd1718:BCD_Out <= 12'b000100000101;
		12'd1719:BCD_Out <= 12'b000100000101;
		12'd1720:BCD_Out <= 12'b000100000101;
		12'd1721:BCD_Out <= 12'b000100000101;
		12'd1722:BCD_Out <= 12'b000100000101;
		12'd1723:BCD_Out <= 12'b000100000101;
		12'd1724:BCD_Out <= 12'b000100000101;
		12'd1725:BCD_Out <= 12'b000100000101;
		12'd1726:BCD_Out <= 12'b000100000101;
		12'd1727:BCD_Out <= 12'b000100000101;
		12'd1728:BCD_Out <= 12'b000100000101;
		12'd1729:BCD_Out <= 12'b000100000110;
		12'd1730:BCD_Out <= 12'b000100000110;
		12'd1731:BCD_Out <= 12'b000100000110;
		12'd1732:BCD_Out <= 12'b000100000110;
		12'd1733:BCD_Out <= 12'b000100000110;
		12'd1734:BCD_Out <= 12'b000100000110;
		12'd1735:BCD_Out <= 12'b000100000110;
		12'd1736:BCD_Out <= 12'b000100000110;
		12'd1737:BCD_Out <= 12'b000100000110;
		12'd1738:BCD_Out <= 12'b000100000110;
		12'd1739:BCD_Out <= 12'b000100000110;
		12'd1740:BCD_Out <= 12'b000100000110;
		12'd1741:BCD_Out <= 12'b000100000110;
		12'd1742:BCD_Out <= 12'b000100000110;
		12'd1743:BCD_Out <= 12'b000100000110;
		12'd1744:BCD_Out <= 12'b000100000110;
		12'd1745:BCD_Out <= 12'b000100000111;
		12'd1746:BCD_Out <= 12'b000100000111;
		12'd1747:BCD_Out <= 12'b000100000111;
		12'd1748:BCD_Out <= 12'b000100000111;
		12'd1749:BCD_Out <= 12'b000100000111;
		12'd1750:BCD_Out <= 12'b000100000111;
		12'd1751:BCD_Out <= 12'b000100000111;
		12'd1752:BCD_Out <= 12'b000100000111;
		12'd1753:BCD_Out <= 12'b000100000111;
		12'd1754:BCD_Out <= 12'b000100000111;
		12'd1755:BCD_Out <= 12'b000100000111;
		12'd1756:BCD_Out <= 12'b000100000111;
		12'd1757:BCD_Out <= 12'b000100000111;
		12'd1758:BCD_Out <= 12'b000100000111;
		12'd1759:BCD_Out <= 12'b000100000111;
		12'd1760:BCD_Out <= 12'b000100000111;
		12'd1761:BCD_Out <= 12'b000100001000;
		12'd1762:BCD_Out <= 12'b000100001000;
		12'd1763:BCD_Out <= 12'b000100001000;
		12'd1764:BCD_Out <= 12'b000100001000;
		12'd1765:BCD_Out <= 12'b000100001000;
		12'd1766:BCD_Out <= 12'b000100001000;
		12'd1767:BCD_Out <= 12'b000100001000;
		12'd1768:BCD_Out <= 12'b000100001000;
		12'd1769:BCD_Out <= 12'b000100001000;
		12'd1770:BCD_Out <= 12'b000100001000;
		12'd1771:BCD_Out <= 12'b000100001000;
		12'd1772:BCD_Out <= 12'b000100001000;
		12'd1773:BCD_Out <= 12'b000100001000;
		12'd1774:BCD_Out <= 12'b000100001000;
		12'd1775:BCD_Out <= 12'b000100001000;
		12'd1776:BCD_Out <= 12'b000100001000;
		12'd1777:BCD_Out <= 12'b000100001000;
		12'd1778:BCD_Out <= 12'b000100001001;
		12'd1779:BCD_Out <= 12'b000100001001;
		12'd1780:BCD_Out <= 12'b000100001001;
		12'd1781:BCD_Out <= 12'b000100001001;
		12'd1782:BCD_Out <= 12'b000100001001;
		12'd1783:BCD_Out <= 12'b000100001001;
		12'd1784:BCD_Out <= 12'b000100001001;
		12'd1785:BCD_Out <= 12'b000100001001;
		12'd1786:BCD_Out <= 12'b000100001001;
		12'd1787:BCD_Out <= 12'b000100001001;
		12'd1788:BCD_Out <= 12'b000100001001;
		12'd1789:BCD_Out <= 12'b000100001001;
		12'd1790:BCD_Out <= 12'b000100001001;
		12'd1791:BCD_Out <= 12'b000100001001;
		12'd1792:BCD_Out <= 12'b000100001001;
		12'd1793:BCD_Out <= 12'b000100001001;
		12'd1794:BCD_Out <= 12'b000100010000;
		12'd1795:BCD_Out <= 12'b000100010000;
		12'd1796:BCD_Out <= 12'b000100010000;
		12'd1797:BCD_Out <= 12'b000100010000;
		12'd1798:BCD_Out <= 12'b000100010000;
		12'd1799:BCD_Out <= 12'b000100010000;
		12'd1800:BCD_Out <= 12'b000100010000;
		12'd1801:BCD_Out <= 12'b000100010000;
		12'd1802:BCD_Out <= 12'b000100010000;
		12'd1803:BCD_Out <= 12'b000100010000;
		12'd1804:BCD_Out <= 12'b000100010000;
		12'd1805:BCD_Out <= 12'b000100010000;
		12'd1806:BCD_Out <= 12'b000100010000;
		12'd1807:BCD_Out <= 12'b000100010000;
		12'd1808:BCD_Out <= 12'b000100010000;
		12'd1809:BCD_Out <= 12'b000100010000;
		12'd1810:BCD_Out <= 12'b000100010001;
		12'd1811:BCD_Out <= 12'b000100010001;
		12'd1812:BCD_Out <= 12'b000100010001;
		12'd1813:BCD_Out <= 12'b000100010001;
		12'd1814:BCD_Out <= 12'b000100010001;
		12'd1815:BCD_Out <= 12'b000100010001;
		12'd1816:BCD_Out <= 12'b000100010001;
		12'd1817:BCD_Out <= 12'b000100010001;
		12'd1818:BCD_Out <= 12'b000100010001;
		12'd1819:BCD_Out <= 12'b000100010001;
		12'd1820:BCD_Out <= 12'b000100010001;
		12'd1821:BCD_Out <= 12'b000100010001;
		12'd1822:BCD_Out <= 12'b000100010001;
		12'd1823:BCD_Out <= 12'b000100010001;
		12'd1824:BCD_Out <= 12'b000100010001;
		12'd1825:BCD_Out <= 12'b000100010001;
		12'd1826:BCD_Out <= 12'b000100010001;
		12'd1827:BCD_Out <= 12'b000100010010;
		12'd1828:BCD_Out <= 12'b000100010010;
		12'd1829:BCD_Out <= 12'b000100010010;
		12'd1830:BCD_Out <= 12'b000100010010;
		12'd1831:BCD_Out <= 12'b000100010010;
		12'd1832:BCD_Out <= 12'b000100010010;
		12'd1833:BCD_Out <= 12'b000100010010;
		12'd1834:BCD_Out <= 12'b000100010010;
		12'd1835:BCD_Out <= 12'b000100010010;
		12'd1836:BCD_Out <= 12'b000100010010;
		12'd1837:BCD_Out <= 12'b000100010010;
		12'd1838:BCD_Out <= 12'b000100010010;
		12'd1839:BCD_Out <= 12'b000100010010;
		12'd1840:BCD_Out <= 12'b000100010010;
		12'd1841:BCD_Out <= 12'b000100010010;
		12'd1842:BCD_Out <= 12'b000100010010;
		12'd1843:BCD_Out <= 12'b000100010011;
		12'd1844:BCD_Out <= 12'b000100010011;
		12'd1845:BCD_Out <= 12'b000100010011;
		12'd1846:BCD_Out <= 12'b000100010011;
		12'd1847:BCD_Out <= 12'b000100010011;
		12'd1848:BCD_Out <= 12'b000100010011;
		12'd1849:BCD_Out <= 12'b000100010011;
		12'd1850:BCD_Out <= 12'b000100010011;
		12'd1851:BCD_Out <= 12'b000100010011;
		12'd1852:BCD_Out <= 12'b000100010011;
		12'd1853:BCD_Out <= 12'b000100010011;
		12'd1854:BCD_Out <= 12'b000100010011;
		12'd1855:BCD_Out <= 12'b000100010011;
		12'd1856:BCD_Out <= 12'b000100010011;
		12'd1857:BCD_Out <= 12'b000100010011;
		12'd1858:BCD_Out <= 12'b000100010011;
		12'd1859:BCD_Out <= 12'b000100010011;
		12'd1860:BCD_Out <= 12'b000100010100;
		12'd1861:BCD_Out <= 12'b000100010100;
		12'd1862:BCD_Out <= 12'b000100010100;
		12'd1863:BCD_Out <= 12'b000100010100;
		12'd1864:BCD_Out <= 12'b000100010100;
		12'd1865:BCD_Out <= 12'b000100010100;
		12'd1866:BCD_Out <= 12'b000100010100;
		12'd1867:BCD_Out <= 12'b000100010100;
		12'd1868:BCD_Out <= 12'b000100010100;
		12'd1869:BCD_Out <= 12'b000100010100;
		12'd1870:BCD_Out <= 12'b000100010100;
		12'd1871:BCD_Out <= 12'b000100010100;
		12'd1872:BCD_Out <= 12'b000100010100;
		12'd1873:BCD_Out <= 12'b000100010100;
		12'd1874:BCD_Out <= 12'b000100010100;
		12'd1875:BCD_Out <= 12'b000100010100;
		12'd1876:BCD_Out <= 12'b000100010101;
		12'd1877:BCD_Out <= 12'b000100010101;
		12'd1878:BCD_Out <= 12'b000100010101;
		12'd1879:BCD_Out <= 12'b000100010101;
		12'd1880:BCD_Out <= 12'b000100010101;
		12'd1881:BCD_Out <= 12'b000100010101;
		12'd1882:BCD_Out <= 12'b000100010101;
		12'd1883:BCD_Out <= 12'b000100010101;
		12'd1884:BCD_Out <= 12'b000100010101;
		12'd1885:BCD_Out <= 12'b000100010101;
		12'd1886:BCD_Out <= 12'b000100010101;
		12'd1887:BCD_Out <= 12'b000100010101;
		12'd1888:BCD_Out <= 12'b000100010101;
		12'd1889:BCD_Out <= 12'b000100010101;
		12'd1890:BCD_Out <= 12'b000100010101;
		12'd1891:BCD_Out <= 12'b000100010101;
		12'd1892:BCD_Out <= 12'b000100010110;
		12'd1893:BCD_Out <= 12'b000100010110;
		12'd1894:BCD_Out <= 12'b000100010110;
		12'd1895:BCD_Out <= 12'b000100010110;
		12'd1896:BCD_Out <= 12'b000100010110;
		12'd1897:BCD_Out <= 12'b000100010110;
		12'd1898:BCD_Out <= 12'b000100010110;
		12'd1899:BCD_Out <= 12'b000100010110;
		12'd1900:BCD_Out <= 12'b000100010110;
		12'd1901:BCD_Out <= 12'b000100010110;
		12'd1902:BCD_Out <= 12'b000100010110;
		12'd1903:BCD_Out <= 12'b000100010110;
		12'd1904:BCD_Out <= 12'b000100010110;
		12'd1905:BCD_Out <= 12'b000100010110;
		12'd1906:BCD_Out <= 12'b000100010110;
		12'd1907:BCD_Out <= 12'b000100010110;
		12'd1908:BCD_Out <= 12'b000100010110;
		12'd1909:BCD_Out <= 12'b000100010111;
		12'd1910:BCD_Out <= 12'b000100010111;
		12'd1911:BCD_Out <= 12'b000100010111;
		12'd1912:BCD_Out <= 12'b000100010111;
		12'd1913:BCD_Out <= 12'b000100010111;
		12'd1914:BCD_Out <= 12'b000100010111;
		12'd1915:BCD_Out <= 12'b000100010111;
		12'd1916:BCD_Out <= 12'b000100010111;
		12'd1917:BCD_Out <= 12'b000100010111;
		12'd1918:BCD_Out <= 12'b000100010111;
		12'd1919:BCD_Out <= 12'b000100010111;
		12'd1920:BCD_Out <= 12'b000100010111;
		12'd1921:BCD_Out <= 12'b000100010111;
		12'd1922:BCD_Out <= 12'b000100010111;
		12'd1923:BCD_Out <= 12'b000100010111;
		12'd1924:BCD_Out <= 12'b000100010111;
		12'd1925:BCD_Out <= 12'b000100011000;
		12'd1926:BCD_Out <= 12'b000100011000;
		12'd1927:BCD_Out <= 12'b000100011000;
		12'd1928:BCD_Out <= 12'b000100011000;
		12'd1929:BCD_Out <= 12'b000100011000;
		12'd1930:BCD_Out <= 12'b000100011000;
		12'd1931:BCD_Out <= 12'b000100011000;
		12'd1932:BCD_Out <= 12'b000100011000;
		12'd1933:BCD_Out <= 12'b000100011000;
		12'd1934:BCD_Out <= 12'b000100011000;
		12'd1935:BCD_Out <= 12'b000100011000;
		12'd1936:BCD_Out <= 12'b000100011000;
		12'd1937:BCD_Out <= 12'b000100011000;
		12'd1938:BCD_Out <= 12'b000100011000;
		12'd1939:BCD_Out <= 12'b000100011000;
		12'd1940:BCD_Out <= 12'b000100011000;
		12'd1941:BCD_Out <= 12'b000100011000;
		12'd1942:BCD_Out <= 12'b000100011001;
		12'd1943:BCD_Out <= 12'b000100011001;
		12'd1944:BCD_Out <= 12'b000100011001;
		12'd1945:BCD_Out <= 12'b000100011001;
		12'd1946:BCD_Out <= 12'b000100011001;
		12'd1947:BCD_Out <= 12'b000100011001;
		12'd1948:BCD_Out <= 12'b000100011001;
		12'd1949:BCD_Out <= 12'b000100011001;
		12'd1950:BCD_Out <= 12'b000100011001;
		12'd1951:BCD_Out <= 12'b000100011001;
		12'd1952:BCD_Out <= 12'b000100011001;
		12'd1953:BCD_Out <= 12'b000100011001;
		12'd1954:BCD_Out <= 12'b000100011001;
		12'd1955:BCD_Out <= 12'b000100011001;
		12'd1956:BCD_Out <= 12'b000100011001;
		12'd1957:BCD_Out <= 12'b000100011001;
		12'd1958:BCD_Out <= 12'b000100100000;
		12'd1959:BCD_Out <= 12'b000100100000;
		12'd1960:BCD_Out <= 12'b000100100000;
		12'd1961:BCD_Out <= 12'b000100100000;
		12'd1962:BCD_Out <= 12'b000100100000;
		12'd1963:BCD_Out <= 12'b000100100000;
		12'd1964:BCD_Out <= 12'b000100100000;
		12'd1965:BCD_Out <= 12'b000100100000;
		12'd1966:BCD_Out <= 12'b000100100000;
		12'd1967:BCD_Out <= 12'b000100100000;
		12'd1968:BCD_Out <= 12'b000100100000;
		12'd1969:BCD_Out <= 12'b000100100000;
		12'd1970:BCD_Out <= 12'b000100100000;
		12'd1971:BCD_Out <= 12'b000100100000;
		12'd1972:BCD_Out <= 12'b000100100000;
		12'd1973:BCD_Out <= 12'b000100100000;
		12'd1974:BCD_Out <= 12'b000100100001;
		12'd1975:BCD_Out <= 12'b000100100001;
		12'd1976:BCD_Out <= 12'b000100100001;
		12'd1977:BCD_Out <= 12'b000100100001;
		12'd1978:BCD_Out <= 12'b000100100001;
		12'd1979:BCD_Out <= 12'b000100100001;
		12'd1980:BCD_Out <= 12'b000100100001;
		12'd1981:BCD_Out <= 12'b000100100001;
		12'd1982:BCD_Out <= 12'b000100100001;
		12'd1983:BCD_Out <= 12'b000100100001;
		12'd1984:BCD_Out <= 12'b000100100001;
		12'd1985:BCD_Out <= 12'b000100100001;
		12'd1986:BCD_Out <= 12'b000100100001;
		12'd1987:BCD_Out <= 12'b000100100001;
		12'd1988:BCD_Out <= 12'b000100100001;
		12'd1989:BCD_Out <= 12'b000100100001;
		12'd1990:BCD_Out <= 12'b000100100001;
		12'd1991:BCD_Out <= 12'b000100100010;
		12'd1992:BCD_Out <= 12'b000100100010;
		12'd1993:BCD_Out <= 12'b000100100010;
		12'd1994:BCD_Out <= 12'b000100100010;
		12'd1995:BCD_Out <= 12'b000100100010;
		12'd1996:BCD_Out <= 12'b000100100010;
		12'd1997:BCD_Out <= 12'b000100100010;
		12'd1998:BCD_Out <= 12'b000100100010;
		12'd1999:BCD_Out <= 12'b000100100010;
		12'd2000:BCD_Out <= 12'b000100100010;
		12'd2001:BCD_Out <= 12'b000100100010;
		12'd2002:BCD_Out <= 12'b000100100010;
		12'd2003:BCD_Out <= 12'b000100100010;
		12'd2004:BCD_Out <= 12'b000100100010;
		12'd2005:BCD_Out <= 12'b000100100010;
		12'd2006:BCD_Out <= 12'b000100100010;
		12'd2007:BCD_Out <= 12'b000100100011;
		12'd2008:BCD_Out <= 12'b000100100011;
		12'd2009:BCD_Out <= 12'b000100100011;
		12'd2010:BCD_Out <= 12'b000100100011;
		12'd2011:BCD_Out <= 12'b000100100011;
		12'd2012:BCD_Out <= 12'b000100100011;
		12'd2013:BCD_Out <= 12'b000100100011;
		12'd2014:BCD_Out <= 12'b000100100011;
		12'd2015:BCD_Out <= 12'b000100100011;
		12'd2016:BCD_Out <= 12'b000100100011;
		12'd2017:BCD_Out <= 12'b000100100011;
		12'd2018:BCD_Out <= 12'b000100100011;
		12'd2019:BCD_Out <= 12'b000100100011;
		12'd2020:BCD_Out <= 12'b000100100011;
		12'd2021:BCD_Out <= 12'b000100100011;
		12'd2022:BCD_Out <= 12'b000100100011;
		12'd2023:BCD_Out <= 12'b000100100100;
		12'd2024:BCD_Out <= 12'b000100100100;
		12'd2025:BCD_Out <= 12'b000100100100;
		12'd2026:BCD_Out <= 12'b000100100100;
		12'd2027:BCD_Out <= 12'b000100100100;
		12'd2028:BCD_Out <= 12'b000100100100;
		12'd2029:BCD_Out <= 12'b000100100100;
		12'd2030:BCD_Out <= 12'b000100100100;
		12'd2031:BCD_Out <= 12'b000100100100;
		12'd2032:BCD_Out <= 12'b000100100100;
		12'd2033:BCD_Out <= 12'b000100100100;
		12'd2034:BCD_Out <= 12'b000100100100;
		12'd2035:BCD_Out <= 12'b000100100100;
		12'd2036:BCD_Out <= 12'b000100100100;
		12'd2037:BCD_Out <= 12'b000100100100;
		12'd2038:BCD_Out <= 12'b000100100100;
		12'd2039:BCD_Out <= 12'b000100100100;
		12'd2040:BCD_Out <= 12'b000100100101;
		12'd2041:BCD_Out <= 12'b000100100101;
		12'd2042:BCD_Out <= 12'b000100100101;
		12'd2043:BCD_Out <= 12'b000100100101;
		12'd2044:BCD_Out <= 12'b000100100101;
		12'd2045:BCD_Out <= 12'b000100100101;
		12'd2046:BCD_Out <= 12'b000100100101;
		12'd2047:BCD_Out <= 12'b000100100101;
		12'd2048:BCD_Out <= 12'b000100100101;
		12'd2049:BCD_Out <= 12'b000100100101;
		12'd2050:BCD_Out <= 12'b000100100101;
		12'd2051:BCD_Out <= 12'b000100100101;
		12'd2052:BCD_Out <= 12'b000100100101;
		12'd2053:BCD_Out <= 12'b000100100101;
		12'd2054:BCD_Out <= 12'b000100100101;
		12'd2055:BCD_Out <= 12'b000100100101;
		12'd2056:BCD_Out <= 12'b000100100110;
		12'd2057:BCD_Out <= 12'b000100100110;
		12'd2058:BCD_Out <= 12'b000100100110;
		12'd2059:BCD_Out <= 12'b000100100110;
		12'd2060:BCD_Out <= 12'b000100100110;
		12'd2061:BCD_Out <= 12'b000100100110;
		12'd2062:BCD_Out <= 12'b000100100110;
		12'd2063:BCD_Out <= 12'b000100100110;
		12'd2064:BCD_Out <= 12'b000100100110;
		12'd2065:BCD_Out <= 12'b000100100110;
		12'd2066:BCD_Out <= 12'b000100100110;
		12'd2067:BCD_Out <= 12'b000100100110;
		12'd2068:BCD_Out <= 12'b000100100110;
		12'd2069:BCD_Out <= 12'b000100100110;
		12'd2070:BCD_Out <= 12'b000100100110;
		12'd2071:BCD_Out <= 12'b000100100110;
		12'd2072:BCD_Out <= 12'b000100100110;
		12'd2073:BCD_Out <= 12'b000100100111;
		12'd2074:BCD_Out <= 12'b000100100111;
		12'd2075:BCD_Out <= 12'b000100100111;
		12'd2076:BCD_Out <= 12'b000100100111;
		12'd2077:BCD_Out <= 12'b000100100111;
		12'd2078:BCD_Out <= 12'b000100100111;
		12'd2079:BCD_Out <= 12'b000100100111;
		12'd2080:BCD_Out <= 12'b000100100111;
		12'd2081:BCD_Out <= 12'b000100100111;
		12'd2082:BCD_Out <= 12'b000100100111;
		12'd2083:BCD_Out <= 12'b000100100111;
		12'd2084:BCD_Out <= 12'b000100100111;
		12'd2085:BCD_Out <= 12'b000100100111;
		12'd2086:BCD_Out <= 12'b000100100111;
		12'd2087:BCD_Out <= 12'b000100100111;
		12'd2088:BCD_Out <= 12'b000100100111;
		12'd2089:BCD_Out <= 12'b000100101000;
		12'd2090:BCD_Out <= 12'b000100101000;
		12'd2091:BCD_Out <= 12'b000100101000;
		12'd2092:BCD_Out <= 12'b000100101000;
		12'd2093:BCD_Out <= 12'b000100101000;
		12'd2094:BCD_Out <= 12'b000100101000;
		12'd2095:BCD_Out <= 12'b000100101000;
		12'd2096:BCD_Out <= 12'b000100101000;
		12'd2097:BCD_Out <= 12'b000100101000;
		12'd2098:BCD_Out <= 12'b000100101000;
		12'd2099:BCD_Out <= 12'b000100101000;
		12'd2100:BCD_Out <= 12'b000100101000;
		12'd2101:BCD_Out <= 12'b000100101000;
		12'd2102:BCD_Out <= 12'b000100101000;
		12'd2103:BCD_Out <= 12'b000100101000;
		12'd2104:BCD_Out <= 12'b000100101000;
		12'd2105:BCD_Out <= 12'b000100101001;
		12'd2106:BCD_Out <= 12'b000100101001;
		12'd2107:BCD_Out <= 12'b000100101001;
		12'd2108:BCD_Out <= 12'b000100101001;
		12'd2109:BCD_Out <= 12'b000100101001;
		12'd2110:BCD_Out <= 12'b000100101001;
		12'd2111:BCD_Out <= 12'b000100101001;
		12'd2112:BCD_Out <= 12'b000100101001;
		12'd2113:BCD_Out <= 12'b000100101001;
		12'd2114:BCD_Out <= 12'b000100101001;
		12'd2115:BCD_Out <= 12'b000100101001;
		12'd2116:BCD_Out <= 12'b000100101001;
		12'd2117:BCD_Out <= 12'b000100101001;
		12'd2118:BCD_Out <= 12'b000100101001;
		12'd2119:BCD_Out <= 12'b000100101001;
		12'd2120:BCD_Out <= 12'b000100101001;
		12'd2121:BCD_Out <= 12'b000100101001;
		12'd2122:BCD_Out <= 12'b000100110000;
		12'd2123:BCD_Out <= 12'b000100110000;
		12'd2124:BCD_Out <= 12'b000100110000;
		12'd2125:BCD_Out <= 12'b000100110000;
		12'd2126:BCD_Out <= 12'b000100110000;
		12'd2127:BCD_Out <= 12'b000100110000;
		12'd2128:BCD_Out <= 12'b000100110000;
		12'd2129:BCD_Out <= 12'b000100110000;
		12'd2130:BCD_Out <= 12'b000100110000;
		12'd2131:BCD_Out <= 12'b000100110000;
		12'd2132:BCD_Out <= 12'b000100110000;
		12'd2133:BCD_Out <= 12'b000100110000;
		12'd2134:BCD_Out <= 12'b000100110000;
		12'd2135:BCD_Out <= 12'b000100110000;
		12'd2136:BCD_Out <= 12'b000100110000;
		12'd2137:BCD_Out <= 12'b000100110000;
		12'd2138:BCD_Out <= 12'b000100110001;
		12'd2139:BCD_Out <= 12'b000100110001;
		12'd2140:BCD_Out <= 12'b000100110001;
		12'd2141:BCD_Out <= 12'b000100110001;
		12'd2142:BCD_Out <= 12'b000100110001;
		12'd2143:BCD_Out <= 12'b000100110001;
		12'd2144:BCD_Out <= 12'b000100110001;
		12'd2145:BCD_Out <= 12'b000100110001;
		12'd2146:BCD_Out <= 12'b000100110001;
		12'd2147:BCD_Out <= 12'b000100110001;
		12'd2148:BCD_Out <= 12'b000100110001;
		12'd2149:BCD_Out <= 12'b000100110001;
		12'd2150:BCD_Out <= 12'b000100110001;
		12'd2151:BCD_Out <= 12'b000100110001;
		12'd2152:BCD_Out <= 12'b000100110001;
		12'd2153:BCD_Out <= 12'b000100110001;
		12'd2154:BCD_Out <= 12'b000100110010;
		12'd2155:BCD_Out <= 12'b000100110010;
		12'd2156:BCD_Out <= 12'b000100110010;
		12'd2157:BCD_Out <= 12'b000100110010;
		12'd2158:BCD_Out <= 12'b000100110010;
		12'd2159:BCD_Out <= 12'b000100110010;
		12'd2160:BCD_Out <= 12'b000100110010;
		12'd2161:BCD_Out <= 12'b000100110010;
		12'd2162:BCD_Out <= 12'b000100110010;
		12'd2163:BCD_Out <= 12'b000100110010;
		12'd2164:BCD_Out <= 12'b000100110010;
		12'd2165:BCD_Out <= 12'b000100110010;
		12'd2166:BCD_Out <= 12'b000100110010;
		12'd2167:BCD_Out <= 12'b000100110010;
		12'd2168:BCD_Out <= 12'b000100110010;
		12'd2169:BCD_Out <= 12'b000100110010;
		12'd2170:BCD_Out <= 12'b000100110010;
		12'd2171:BCD_Out <= 12'b000100110011;
		12'd2172:BCD_Out <= 12'b000100110011;
		12'd2173:BCD_Out <= 12'b000100110011;
		12'd2174:BCD_Out <= 12'b000100110011;
		12'd2175:BCD_Out <= 12'b000100110011;
		12'd2176:BCD_Out <= 12'b000100110011;
		12'd2177:BCD_Out <= 12'b000100110011;
		12'd2178:BCD_Out <= 12'b000100110011;
		12'd2179:BCD_Out <= 12'b000100110011;
		12'd2180:BCD_Out <= 12'b000100110011;
		12'd2181:BCD_Out <= 12'b000100110011;
		12'd2182:BCD_Out <= 12'b000100110011;
		12'd2183:BCD_Out <= 12'b000100110011;
		12'd2184:BCD_Out <= 12'b000100110011;
		12'd2185:BCD_Out <= 12'b000100110011;
		12'd2186:BCD_Out <= 12'b000100110011;
		12'd2187:BCD_Out <= 12'b000100110100;
		12'd2188:BCD_Out <= 12'b000100110100;
		12'd2189:BCD_Out <= 12'b000100110100;
		12'd2190:BCD_Out <= 12'b000100110100;
		12'd2191:BCD_Out <= 12'b000100110100;
		12'd2192:BCD_Out <= 12'b000100110100;
		12'd2193:BCD_Out <= 12'b000100110100;
		12'd2194:BCD_Out <= 12'b000100110100;
		12'd2195:BCD_Out <= 12'b000100110100;
		12'd2196:BCD_Out <= 12'b000100110100;
		12'd2197:BCD_Out <= 12'b000100110100;
		12'd2198:BCD_Out <= 12'b000100110100;
		12'd2199:BCD_Out <= 12'b000100110100;
		12'd2200:BCD_Out <= 12'b000100110100;
		12'd2201:BCD_Out <= 12'b000100110100;
		12'd2202:BCD_Out <= 12'b000100110100;
		12'd2203:BCD_Out <= 12'b000100110100;
		12'd2204:BCD_Out <= 12'b000100110101;
		12'd2205:BCD_Out <= 12'b000100110101;
		12'd2206:BCD_Out <= 12'b000100110101;
		12'd2207:BCD_Out <= 12'b000100110101;
		12'd2208:BCD_Out <= 12'b000100110101;
		12'd2209:BCD_Out <= 12'b000100110101;
		12'd2210:BCD_Out <= 12'b000100110101;
		12'd2211:BCD_Out <= 12'b000100110101;
		12'd2212:BCD_Out <= 12'b000100110101;
		12'd2213:BCD_Out <= 12'b000100110101;
		12'd2214:BCD_Out <= 12'b000100110101;
		12'd2215:BCD_Out <= 12'b000100110101;
		12'd2216:BCD_Out <= 12'b000100110101;
		12'd2217:BCD_Out <= 12'b000100110101;
		12'd2218:BCD_Out <= 12'b000100110101;
		12'd2219:BCD_Out <= 12'b000100110101;
		12'd2220:BCD_Out <= 12'b000100110110;
		12'd2221:BCD_Out <= 12'b000100110110;
		12'd2222:BCD_Out <= 12'b000100110110;
		12'd2223:BCD_Out <= 12'b000100110110;
		12'd2224:BCD_Out <= 12'b000100110110;
		12'd2225:BCD_Out <= 12'b000100110110;
		12'd2226:BCD_Out <= 12'b000100110110;
		12'd2227:BCD_Out <= 12'b000100110110;
		12'd2228:BCD_Out <= 12'b000100110110;
		12'd2229:BCD_Out <= 12'b000100110110;
		12'd2230:BCD_Out <= 12'b000100110110;
		12'd2231:BCD_Out <= 12'b000100110110;
		12'd2232:BCD_Out <= 12'b000100110110;
		12'd2233:BCD_Out <= 12'b000100110110;
		12'd2234:BCD_Out <= 12'b000100110110;
		12'd2235:BCD_Out <= 12'b000100110110;
		12'd2236:BCD_Out <= 12'b000100110111;
		12'd2237:BCD_Out <= 12'b000100110111;
		12'd2238:BCD_Out <= 12'b000100110111;
		12'd2239:BCD_Out <= 12'b000100110111;
		12'd2240:BCD_Out <= 12'b000100110111;
		12'd2241:BCD_Out <= 12'b000100110111;
		12'd2242:BCD_Out <= 12'b000100110111;
		12'd2243:BCD_Out <= 12'b000100110111;
		12'd2244:BCD_Out <= 12'b000100110111;
		12'd2245:BCD_Out <= 12'b000100110111;
		12'd2246:BCD_Out <= 12'b000100110111;
		12'd2247:BCD_Out <= 12'b000100110111;
		12'd2248:BCD_Out <= 12'b000100110111;
		12'd2249:BCD_Out <= 12'b000100110111;
		12'd2250:BCD_Out <= 12'b000100110111;
		12'd2251:BCD_Out <= 12'b000100110111;
		12'd2252:BCD_Out <= 12'b000100110111;
		12'd2253:BCD_Out <= 12'b000100111000;
		12'd2254:BCD_Out <= 12'b000100111000;
		12'd2255:BCD_Out <= 12'b000100111000;
		12'd2256:BCD_Out <= 12'b000100111000;
		12'd2257:BCD_Out <= 12'b000100111000;
		12'd2258:BCD_Out <= 12'b000100111000;
		12'd2259:BCD_Out <= 12'b000100111000;
		12'd2260:BCD_Out <= 12'b000100111000;
		12'd2261:BCD_Out <= 12'b000100111000;
		12'd2262:BCD_Out <= 12'b000100111000;
		12'd2263:BCD_Out <= 12'b000100111000;
		12'd2264:BCD_Out <= 12'b000100111000;
		12'd2265:BCD_Out <= 12'b000100111000;
		12'd2266:BCD_Out <= 12'b000100111000;
		12'd2267:BCD_Out <= 12'b000100111000;
		12'd2268:BCD_Out <= 12'b000100111000;
		12'd2269:BCD_Out <= 12'b000100111001;
		12'd2270:BCD_Out <= 12'b000100111001;
		12'd2271:BCD_Out <= 12'b000100111001;
		12'd2272:BCD_Out <= 12'b000100111001;
		12'd2273:BCD_Out <= 12'b000100111001;
		12'd2274:BCD_Out <= 12'b000100111001;
		12'd2275:BCD_Out <= 12'b000100111001;
		12'd2276:BCD_Out <= 12'b000100111001;
		12'd2277:BCD_Out <= 12'b000100111001;
		12'd2278:BCD_Out <= 12'b000100111001;
		12'd2279:BCD_Out <= 12'b000100111001;
		12'd2280:BCD_Out <= 12'b000100111001;
		12'd2281:BCD_Out <= 12'b000100111001;
		12'd2282:BCD_Out <= 12'b000100111001;
		12'd2283:BCD_Out <= 12'b000100111001;
		12'd2284:BCD_Out <= 12'b000100111001;
		12'd2285:BCD_Out <= 12'b000100111001;
		12'd2286:BCD_Out <= 12'b000101000000;
		12'd2287:BCD_Out <= 12'b000101000000;
		12'd2288:BCD_Out <= 12'b000101000000;
		12'd2289:BCD_Out <= 12'b000101000000;
		12'd2290:BCD_Out <= 12'b000101000000;
		12'd2291:BCD_Out <= 12'b000101000000;
		12'd2292:BCD_Out <= 12'b000101000000;
		12'd2293:BCD_Out <= 12'b000101000000;
		12'd2294:BCD_Out <= 12'b000101000000;
		12'd2295:BCD_Out <= 12'b000101000000;
		12'd2296:BCD_Out <= 12'b000101000000;
		12'd2297:BCD_Out <= 12'b000101000000;
		12'd2298:BCD_Out <= 12'b000101000000;
		12'd2299:BCD_Out <= 12'b000101000000;
		12'd2300:BCD_Out <= 12'b000101000000;
		12'd2301:BCD_Out <= 12'b000101000000;
		12'd2302:BCD_Out <= 12'b000101000001;
		12'd2303:BCD_Out <= 12'b000101000001;
		12'd2304:BCD_Out <= 12'b000101000001;
		12'd2305:BCD_Out <= 12'b000101000001;
		12'd2306:BCD_Out <= 12'b000101000001;
		12'd2307:BCD_Out <= 12'b000101000001;
		12'd2308:BCD_Out <= 12'b000101000001;
		12'd2309:BCD_Out <= 12'b000101000001;
		12'd2310:BCD_Out <= 12'b000101000001;
		12'd2311:BCD_Out <= 12'b000101000001;
		12'd2312:BCD_Out <= 12'b000101000001;
		12'd2313:BCD_Out <= 12'b000101000001;
		12'd2314:BCD_Out <= 12'b000101000001;
		12'd2315:BCD_Out <= 12'b000101000001;
		12'd2316:BCD_Out <= 12'b000101000001;
		12'd2317:BCD_Out <= 12'b000101000001;
		12'd2318:BCD_Out <= 12'b000101000010;
		12'd2319:BCD_Out <= 12'b000101000010;
		12'd2320:BCD_Out <= 12'b000101000010;
		12'd2321:BCD_Out <= 12'b000101000010;
		12'd2322:BCD_Out <= 12'b000101000010;
		12'd2323:BCD_Out <= 12'b000101000010;
		12'd2324:BCD_Out <= 12'b000101000010;
		12'd2325:BCD_Out <= 12'b000101000010;
		12'd2326:BCD_Out <= 12'b000101000010;
		12'd2327:BCD_Out <= 12'b000101000010;
		12'd2328:BCD_Out <= 12'b000101000010;
		12'd2329:BCD_Out <= 12'b000101000010;
		12'd2330:BCD_Out <= 12'b000101000010;
		12'd2331:BCD_Out <= 12'b000101000010;
		12'd2332:BCD_Out <= 12'b000101000010;
		12'd2333:BCD_Out <= 12'b000101000010;
		12'd2334:BCD_Out <= 12'b000101000010;
		12'd2335:BCD_Out <= 12'b000101000011;
		12'd2336:BCD_Out <= 12'b000101000011;
		12'd2337:BCD_Out <= 12'b000101000011;
		12'd2338:BCD_Out <= 12'b000101000011;
		12'd2339:BCD_Out <= 12'b000101000011;
		12'd2340:BCD_Out <= 12'b000101000011;
		12'd2341:BCD_Out <= 12'b000101000011;
		12'd2342:BCD_Out <= 12'b000101000011;
		12'd2343:BCD_Out <= 12'b000101000011;
		12'd2344:BCD_Out <= 12'b000101000011;
		12'd2345:BCD_Out <= 12'b000101000011;
		12'd2346:BCD_Out <= 12'b000101000011;
		12'd2347:BCD_Out <= 12'b000101000011;
		12'd2348:BCD_Out <= 12'b000101000011;
		12'd2349:BCD_Out <= 12'b000101000011;
		12'd2350:BCD_Out <= 12'b000101000011;
		12'd2351:BCD_Out <= 12'b000101000100;
		12'd2352:BCD_Out <= 12'b000101000100;
		12'd2353:BCD_Out <= 12'b000101000100;
		12'd2354:BCD_Out <= 12'b000101000100;
		12'd2355:BCD_Out <= 12'b000101000100;
		12'd2356:BCD_Out <= 12'b000101000100;
		12'd2357:BCD_Out <= 12'b000101000100;
		12'd2358:BCD_Out <= 12'b000101000100;
		12'd2359:BCD_Out <= 12'b000101000100;
		12'd2360:BCD_Out <= 12'b000101000100;
		12'd2361:BCD_Out <= 12'b000101000100;
		12'd2362:BCD_Out <= 12'b000101000100;
		12'd2363:BCD_Out <= 12'b000101000100;
		12'd2364:BCD_Out <= 12'b000101000100;
		12'd2365:BCD_Out <= 12'b000101000100;
		12'd2366:BCD_Out <= 12'b000101000100;
		12'd2367:BCD_Out <= 12'b000101000101;
		12'd2368:BCD_Out <= 12'b000101000101;
		12'd2369:BCD_Out <= 12'b000101000101;
		12'd2370:BCD_Out <= 12'b000101000101;
		12'd2371:BCD_Out <= 12'b000101000101;
		12'd2372:BCD_Out <= 12'b000101000101;
		12'd2373:BCD_Out <= 12'b000101000101;
		12'd2374:BCD_Out <= 12'b000101000101;
		12'd2375:BCD_Out <= 12'b000101000101;
		12'd2376:BCD_Out <= 12'b000101000101;
		12'd2377:BCD_Out <= 12'b000101000101;
		12'd2378:BCD_Out <= 12'b000101000101;
		12'd2379:BCD_Out <= 12'b000101000101;
		12'd2380:BCD_Out <= 12'b000101000101;
		12'd2381:BCD_Out <= 12'b000101000101;
		12'd2382:BCD_Out <= 12'b000101000101;
		12'd2383:BCD_Out <= 12'b000101000101;
		12'd2384:BCD_Out <= 12'b000101000110;
		12'd2385:BCD_Out <= 12'b000101000110;
		12'd2386:BCD_Out <= 12'b000101000110;
		12'd2387:BCD_Out <= 12'b000101000110;
		12'd2388:BCD_Out <= 12'b000101000110;
		12'd2389:BCD_Out <= 12'b000101000110;
		12'd2390:BCD_Out <= 12'b000101000110;
		12'd2391:BCD_Out <= 12'b000101000110;
		12'd2392:BCD_Out <= 12'b000101000110;
		12'd2393:BCD_Out <= 12'b000101000110;
		12'd2394:BCD_Out <= 12'b000101000110;
		12'd2395:BCD_Out <= 12'b000101000110;
		12'd2396:BCD_Out <= 12'b000101000110;
		12'd2397:BCD_Out <= 12'b000101000110;
		12'd2398:BCD_Out <= 12'b000101000110;
		12'd2399:BCD_Out <= 12'b000101000110;
		12'd2400:BCD_Out <= 12'b000101000111;
		12'd2401:BCD_Out <= 12'b000101000111;
		12'd2402:BCD_Out <= 12'b000101000111;
		12'd2403:BCD_Out <= 12'b000101000111;
		12'd2404:BCD_Out <= 12'b000101000111;
		12'd2405:BCD_Out <= 12'b000101000111;
		12'd2406:BCD_Out <= 12'b000101000111;
		12'd2407:BCD_Out <= 12'b000101000111;
		12'd2408:BCD_Out <= 12'b000101000111;
		12'd2409:BCD_Out <= 12'b000101000111;
		12'd2410:BCD_Out <= 12'b000101000111;
		12'd2411:BCD_Out <= 12'b000101000111;
		12'd2412:BCD_Out <= 12'b000101000111;
		12'd2413:BCD_Out <= 12'b000101000111;
		12'd2414:BCD_Out <= 12'b000101000111;
		12'd2415:BCD_Out <= 12'b000101000111;
		12'd2416:BCD_Out <= 12'b000101000111;
		12'd2417:BCD_Out <= 12'b000101001000;
		12'd2418:BCD_Out <= 12'b000101001000;
		12'd2419:BCD_Out <= 12'b000101001000;
		12'd2420:BCD_Out <= 12'b000101001000;
		12'd2421:BCD_Out <= 12'b000101001000;
		12'd2422:BCD_Out <= 12'b000101001000;
		12'd2423:BCD_Out <= 12'b000101001000;
		12'd2424:BCD_Out <= 12'b000101001000;
		12'd2425:BCD_Out <= 12'b000101001000;
		12'd2426:BCD_Out <= 12'b000101001000;
		12'd2427:BCD_Out <= 12'b000101001000;
		12'd2428:BCD_Out <= 12'b000101001000;
		12'd2429:BCD_Out <= 12'b000101001000;
		12'd2430:BCD_Out <= 12'b000101001000;
		12'd2431:BCD_Out <= 12'b000101001000;
		12'd2432:BCD_Out <= 12'b000101001000;
		12'd2433:BCD_Out <= 12'b000101001001;
		12'd2434:BCD_Out <= 12'b000101001001;
		12'd2435:BCD_Out <= 12'b000101001001;
		12'd2436:BCD_Out <= 12'b000101001001;
		12'd2437:BCD_Out <= 12'b000101001001;
		12'd2438:BCD_Out <= 12'b000101001001;
		12'd2439:BCD_Out <= 12'b000101001001;
		12'd2440:BCD_Out <= 12'b000101001001;
		12'd2441:BCD_Out <= 12'b000101001001;
		12'd2442:BCD_Out <= 12'b000101001001;
		12'd2443:BCD_Out <= 12'b000101001001;
		12'd2444:BCD_Out <= 12'b000101001001;
		12'd2445:BCD_Out <= 12'b000101001001;
		12'd2446:BCD_Out <= 12'b000101001001;
		12'd2447:BCD_Out <= 12'b000101001001;
		12'd2448:BCD_Out <= 12'b000101001001;
		12'd2449:BCD_Out <= 12'b000101010000;
		12'd2450:BCD_Out <= 12'b000101010000;
		12'd2451:BCD_Out <= 12'b000101010000;
		12'd2452:BCD_Out <= 12'b000101010000;
		12'd2453:BCD_Out <= 12'b000101010000;
		12'd2454:BCD_Out <= 12'b000101010000;
		12'd2455:BCD_Out <= 12'b000101010000;
		12'd2456:BCD_Out <= 12'b000101010000;
		12'd2457:BCD_Out <= 12'b000101010000;
		12'd2458:BCD_Out <= 12'b000101010000;
		12'd2459:BCD_Out <= 12'b000101010000;
		12'd2460:BCD_Out <= 12'b000101010000;
		12'd2461:BCD_Out <= 12'b000101010000;
		12'd2462:BCD_Out <= 12'b000101010000;
		12'd2463:BCD_Out <= 12'b000101010000;
		12'd2464:BCD_Out <= 12'b000101010000;
		12'd2465:BCD_Out <= 12'b000101010000;
		12'd2466:BCD_Out <= 12'b000101010001;
		12'd2467:BCD_Out <= 12'b000101010001;
		12'd2468:BCD_Out <= 12'b000101010001;
		12'd2469:BCD_Out <= 12'b000101010001;
		12'd2470:BCD_Out <= 12'b000101010001;
		12'd2471:BCD_Out <= 12'b000101010001;
		12'd2472:BCD_Out <= 12'b000101010001;
		12'd2473:BCD_Out <= 12'b000101010001;
		12'd2474:BCD_Out <= 12'b000101010001;
		12'd2475:BCD_Out <= 12'b000101010001;
		12'd2476:BCD_Out <= 12'b000101010001;
		12'd2477:BCD_Out <= 12'b000101010001;
		12'd2478:BCD_Out <= 12'b000101010001;
		12'd2479:BCD_Out <= 12'b000101010001;
		12'd2480:BCD_Out <= 12'b000101010001;
		12'd2481:BCD_Out <= 12'b000101010001;
		12'd2482:BCD_Out <= 12'b000101010010;
		12'd2483:BCD_Out <= 12'b000101010010;
		12'd2484:BCD_Out <= 12'b000101010010;
		12'd2485:BCD_Out <= 12'b000101010010;
		12'd2486:BCD_Out <= 12'b000101010010;
		12'd2487:BCD_Out <= 12'b000101010010;
		12'd2488:BCD_Out <= 12'b000101010010;
		12'd2489:BCD_Out <= 12'b000101010010;
		12'd2490:BCD_Out <= 12'b000101010010;
		12'd2491:BCD_Out <= 12'b000101010010;
		12'd2492:BCD_Out <= 12'b000101010010;
		12'd2493:BCD_Out <= 12'b000101010010;
		12'd2494:BCD_Out <= 12'b000101010010;
		12'd2495:BCD_Out <= 12'b000101010010;
		12'd2496:BCD_Out <= 12'b000101010010;
		12'd2497:BCD_Out <= 12'b000101010010;
		12'd2498:BCD_Out <= 12'b000101010011;
		12'd2499:BCD_Out <= 12'b000101010011;
		12'd2500:BCD_Out <= 12'b000101010011;
		12'd2501:BCD_Out <= 12'b000101010011;
		12'd2502:BCD_Out <= 12'b000101010011;
		12'd2503:BCD_Out <= 12'b000101010011;
		12'd2504:BCD_Out <= 12'b000101010011;
		12'd2505:BCD_Out <= 12'b000101010011;
		12'd2506:BCD_Out <= 12'b000101010011;
		12'd2507:BCD_Out <= 12'b000101010011;
		12'd2508:BCD_Out <= 12'b000101010011;
		12'd2509:BCD_Out <= 12'b000101010011;
		12'd2510:BCD_Out <= 12'b000101010011;
		12'd2511:BCD_Out <= 12'b000101010011;
		12'd2512:BCD_Out <= 12'b000101010011;
		12'd2513:BCD_Out <= 12'b000101010011;
		12'd2514:BCD_Out <= 12'b000101010011;
		12'd2515:BCD_Out <= 12'b000101010100;
		12'd2516:BCD_Out <= 12'b000101010100;
		12'd2517:BCD_Out <= 12'b000101010100;
		12'd2518:BCD_Out <= 12'b000101010100;
		12'd2519:BCD_Out <= 12'b000101010100;
		12'd2520:BCD_Out <= 12'b000101010100;
		12'd2521:BCD_Out <= 12'b000101010100;
		12'd2522:BCD_Out <= 12'b000101010100;
		12'd2523:BCD_Out <= 12'b000101010100;
		12'd2524:BCD_Out <= 12'b000101010100;
		12'd2525:BCD_Out <= 12'b000101010100;
		12'd2526:BCD_Out <= 12'b000101010100;
		12'd2527:BCD_Out <= 12'b000101010100;
		12'd2528:BCD_Out <= 12'b000101010100;
		12'd2529:BCD_Out <= 12'b000101010100;
		12'd2530:BCD_Out <= 12'b000101010100;
		12'd2531:BCD_Out <= 12'b000101010101;
		12'd2532:BCD_Out <= 12'b000101010101;
		12'd2533:BCD_Out <= 12'b000101010101;
		12'd2534:BCD_Out <= 12'b000101010101;
		12'd2535:BCD_Out <= 12'b000101010101;
		12'd2536:BCD_Out <= 12'b000101010101;
		12'd2537:BCD_Out <= 12'b000101010101;
		12'd2538:BCD_Out <= 12'b000101010101;
		12'd2539:BCD_Out <= 12'b000101010101;
		12'd2540:BCD_Out <= 12'b000101010101;
		12'd2541:BCD_Out <= 12'b000101010101;
		12'd2542:BCD_Out <= 12'b000101010101;
		12'd2543:BCD_Out <= 12'b000101010101;
		12'd2544:BCD_Out <= 12'b000101010101;
		12'd2545:BCD_Out <= 12'b000101010101;
		12'd2546:BCD_Out <= 12'b000101010101;
		12'd2547:BCD_Out <= 12'b000101010101;
		12'd2548:BCD_Out <= 12'b000101010110;
		12'd2549:BCD_Out <= 12'b000101010110;
		12'd2550:BCD_Out <= 12'b000101010110;
		12'd2551:BCD_Out <= 12'b000101010110;
		12'd2552:BCD_Out <= 12'b000101010110;
		12'd2553:BCD_Out <= 12'b000101010110;
		12'd2554:BCD_Out <= 12'b000101010110;
		12'd2555:BCD_Out <= 12'b000101010110;
		12'd2556:BCD_Out <= 12'b000101010110;
		12'd2557:BCD_Out <= 12'b000101010110;
		12'd2558:BCD_Out <= 12'b000101010110;
		12'd2559:BCD_Out <= 12'b000101010110;
		12'd2560:BCD_Out <= 12'b000101010110;
		12'd2561:BCD_Out <= 12'b000101010110;
		12'd2562:BCD_Out <= 12'b000101010110;
		12'd2563:BCD_Out <= 12'b000101010110;
		12'd2564:BCD_Out <= 12'b000101010111;
		12'd2565:BCD_Out <= 12'b000101010111;
		12'd2566:BCD_Out <= 12'b000101010111;
		12'd2567:BCD_Out <= 12'b000101010111;
		12'd2568:BCD_Out <= 12'b000101010111;
		12'd2569:BCD_Out <= 12'b000101010111;
		12'd2570:BCD_Out <= 12'b000101010111;
		12'd2571:BCD_Out <= 12'b000101010111;
		12'd2572:BCD_Out <= 12'b000101010111;
		12'd2573:BCD_Out <= 12'b000101010111;
		12'd2574:BCD_Out <= 12'b000101010111;
		12'd2575:BCD_Out <= 12'b000101010111;
		12'd2576:BCD_Out <= 12'b000101010111;
		12'd2577:BCD_Out <= 12'b000101010111;
		12'd2578:BCD_Out <= 12'b000101010111;
		12'd2579:BCD_Out <= 12'b000101010111;
		12'd2580:BCD_Out <= 12'b000101011000;
		12'd2581:BCD_Out <= 12'b000101011000;
		12'd2582:BCD_Out <= 12'b000101011000;
		12'd2583:BCD_Out <= 12'b000101011000;
		12'd2584:BCD_Out <= 12'b000101011000;
		12'd2585:BCD_Out <= 12'b000101011000;
		12'd2586:BCD_Out <= 12'b000101011000;
		12'd2587:BCD_Out <= 12'b000101011000;
		12'd2588:BCD_Out <= 12'b000101011000;
		12'd2589:BCD_Out <= 12'b000101011000;
		12'd2590:BCD_Out <= 12'b000101011000;
		12'd2591:BCD_Out <= 12'b000101011000;
		12'd2592:BCD_Out <= 12'b000101011000;
		12'd2593:BCD_Out <= 12'b000101011000;
		12'd2594:BCD_Out <= 12'b000101011000;
		12'd2595:BCD_Out <= 12'b000101011000;
		12'd2596:BCD_Out <= 12'b000101011000;
		12'd2597:BCD_Out <= 12'b000101011001;
		12'd2598:BCD_Out <= 12'b000101011001;
		12'd2599:BCD_Out <= 12'b000101011001;
		12'd2600:BCD_Out <= 12'b000101011001;
		12'd2601:BCD_Out <= 12'b000101011001;
		12'd2602:BCD_Out <= 12'b000101011001;
		12'd2603:BCD_Out <= 12'b000101011001;
		12'd2604:BCD_Out <= 12'b000101011001;
		12'd2605:BCD_Out <= 12'b000101011001;
		12'd2606:BCD_Out <= 12'b000101011001;
		12'd2607:BCD_Out <= 12'b000101011001;
		12'd2608:BCD_Out <= 12'b000101011001;
		12'd2609:BCD_Out <= 12'b000101011001;
		12'd2610:BCD_Out <= 12'b000101011001;
		12'd2611:BCD_Out <= 12'b000101011001;
		12'd2612:BCD_Out <= 12'b000101011001;
		12'd2613:BCD_Out <= 12'b000101100000;
		12'd2614:BCD_Out <= 12'b000101100000;
		12'd2615:BCD_Out <= 12'b000101100000;
		12'd2616:BCD_Out <= 12'b000101100000;
		12'd2617:BCD_Out <= 12'b000101100000;
		12'd2618:BCD_Out <= 12'b000101100000;
		12'd2619:BCD_Out <= 12'b000101100000;
		12'd2620:BCD_Out <= 12'b000101100000;
		12'd2621:BCD_Out <= 12'b000101100000;
		12'd2622:BCD_Out <= 12'b000101100000;
		12'd2623:BCD_Out <= 12'b000101100000;
		12'd2624:BCD_Out <= 12'b000101100000;
		12'd2625:BCD_Out <= 12'b000101100000;
		12'd2626:BCD_Out <= 12'b000101100000;
		12'd2627:BCD_Out <= 12'b000101100000;
		12'd2628:BCD_Out <= 12'b000101100000;
		12'd2629:BCD_Out <= 12'b000101100001;
		12'd2630:BCD_Out <= 12'b000101100001;
		12'd2631:BCD_Out <= 12'b000101100001;
		12'd2632:BCD_Out <= 12'b000101100001;
		12'd2633:BCD_Out <= 12'b000101100001;
		12'd2634:BCD_Out <= 12'b000101100001;
		12'd2635:BCD_Out <= 12'b000101100001;
		12'd2636:BCD_Out <= 12'b000101100001;
		12'd2637:BCD_Out <= 12'b000101100001;
		12'd2638:BCD_Out <= 12'b000101100001;
		12'd2639:BCD_Out <= 12'b000101100001;
		12'd2640:BCD_Out <= 12'b000101100001;
		12'd2641:BCD_Out <= 12'b000101100001;
		12'd2642:BCD_Out <= 12'b000101100001;
		12'd2643:BCD_Out <= 12'b000101100001;
		12'd2644:BCD_Out <= 12'b000101100001;
		12'd2645:BCD_Out <= 12'b000101100001;
		12'd2646:BCD_Out <= 12'b000101100010;
		12'd2647:BCD_Out <= 12'b000101100010;
		12'd2648:BCD_Out <= 12'b000101100010;
		12'd2649:BCD_Out <= 12'b000101100010;
		12'd2650:BCD_Out <= 12'b000101100010;
		12'd2651:BCD_Out <= 12'b000101100010;
		12'd2652:BCD_Out <= 12'b000101100010;
		12'd2653:BCD_Out <= 12'b000101100010;
		12'd2654:BCD_Out <= 12'b000101100010;
		12'd2655:BCD_Out <= 12'b000101100010;
		12'd2656:BCD_Out <= 12'b000101100010;
		12'd2657:BCD_Out <= 12'b000101100010;
		12'd2658:BCD_Out <= 12'b000101100010;
		12'd2659:BCD_Out <= 12'b000101100010;
		12'd2660:BCD_Out <= 12'b000101100010;
		12'd2661:BCD_Out <= 12'b000101100010;
		12'd2662:BCD_Out <= 12'b000101100011;
		12'd2663:BCD_Out <= 12'b000101100011;
		12'd2664:BCD_Out <= 12'b000101100011;
		12'd2665:BCD_Out <= 12'b000101100011;
		12'd2666:BCD_Out <= 12'b000101100011;
		12'd2667:BCD_Out <= 12'b000101100011;
		12'd2668:BCD_Out <= 12'b000101100011;
		12'd2669:BCD_Out <= 12'b000101100011;
		12'd2670:BCD_Out <= 12'b000101100011;
		12'd2671:BCD_Out <= 12'b000101100011;
		12'd2672:BCD_Out <= 12'b000101100011;
		12'd2673:BCD_Out <= 12'b000101100011;
		12'd2674:BCD_Out <= 12'b000101100011;
		12'd2675:BCD_Out <= 12'b000101100011;
		12'd2676:BCD_Out <= 12'b000101100011;
		12'd2677:BCD_Out <= 12'b000101100011;
		12'd2678:BCD_Out <= 12'b000101100011;
		12'd2679:BCD_Out <= 12'b000101100100;
		12'd2680:BCD_Out <= 12'b000101100100;
		12'd2681:BCD_Out <= 12'b000101100100;
		12'd2682:BCD_Out <= 12'b000101100100;
		12'd2683:BCD_Out <= 12'b000101100100;
		12'd2684:BCD_Out <= 12'b000101100100;
		12'd2685:BCD_Out <= 12'b000101100100;
		12'd2686:BCD_Out <= 12'b000101100100;
		12'd2687:BCD_Out <= 12'b000101100100;
		12'd2688:BCD_Out <= 12'b000101100100;
		12'd2689:BCD_Out <= 12'b000101100100;
		12'd2690:BCD_Out <= 12'b000101100100;
		12'd2691:BCD_Out <= 12'b000101100100;
		12'd2692:BCD_Out <= 12'b000101100100;
		12'd2693:BCD_Out <= 12'b000101100100;
		12'd2694:BCD_Out <= 12'b000101100100;
		12'd2695:BCD_Out <= 12'b000101100101;
		12'd2696:BCD_Out <= 12'b000101100101;
		12'd2697:BCD_Out <= 12'b000101100101;
		12'd2698:BCD_Out <= 12'b000101100101;
		12'd2699:BCD_Out <= 12'b000101100101;
		12'd2700:BCD_Out <= 12'b000101100101;
		12'd2701:BCD_Out <= 12'b000101100101;
		12'd2702:BCD_Out <= 12'b000101100101;
		12'd2703:BCD_Out <= 12'b000101100101;
		12'd2704:BCD_Out <= 12'b000101100101;
		12'd2705:BCD_Out <= 12'b000101100101;
		12'd2706:BCD_Out <= 12'b000101100101;
		12'd2707:BCD_Out <= 12'b000101100101;
		12'd2708:BCD_Out <= 12'b000101100101;
		12'd2709:BCD_Out <= 12'b000101100101;
		12'd2710:BCD_Out <= 12'b000101100101;
		12'd2711:BCD_Out <= 12'b000101100110;
		12'd2712:BCD_Out <= 12'b000101100110;
		12'd2713:BCD_Out <= 12'b000101100110;
		12'd2714:BCD_Out <= 12'b000101100110;
		12'd2715:BCD_Out <= 12'b000101100110;
		12'd2716:BCD_Out <= 12'b000101100110;
		12'd2717:BCD_Out <= 12'b000101100110;
		12'd2718:BCD_Out <= 12'b000101100110;
		12'd2719:BCD_Out <= 12'b000101100110;
		12'd2720:BCD_Out <= 12'b000101100110;
		12'd2721:BCD_Out <= 12'b000101100110;
		12'd2722:BCD_Out <= 12'b000101100110;
		12'd2723:BCD_Out <= 12'b000101100110;
		12'd2724:BCD_Out <= 12'b000101100110;
		12'd2725:BCD_Out <= 12'b000101100110;
		12'd2726:BCD_Out <= 12'b000101100110;
		12'd2727:BCD_Out <= 12'b000101100110;
		12'd2728:BCD_Out <= 12'b000101100111;
		12'd2729:BCD_Out <= 12'b000101100111;
		12'd2730:BCD_Out <= 12'b000101100111;
		12'd2731:BCD_Out <= 12'b000101100111;
		12'd2732:BCD_Out <= 12'b000101100111;
		12'd2733:BCD_Out <= 12'b000101100111;
		12'd2734:BCD_Out <= 12'b000101100111;
		12'd2735:BCD_Out <= 12'b000101100111;
		12'd2736:BCD_Out <= 12'b000101100111;
		12'd2737:BCD_Out <= 12'b000101100111;
		12'd2738:BCD_Out <= 12'b000101100111;
		12'd2739:BCD_Out <= 12'b000101100111;
		12'd2740:BCD_Out <= 12'b000101100111;
		12'd2741:BCD_Out <= 12'b000101100111;
		12'd2742:BCD_Out <= 12'b000101100111;
		12'd2743:BCD_Out <= 12'b000101100111;
		12'd2744:BCD_Out <= 12'b000101101000;
		12'd2745:BCD_Out <= 12'b000101101000;
		12'd2746:BCD_Out <= 12'b000101101000;
		12'd2747:BCD_Out <= 12'b000101101000;
		12'd2748:BCD_Out <= 12'b000101101000;
		12'd2749:BCD_Out <= 12'b000101101000;
		12'd2750:BCD_Out <= 12'b000101101000;
		12'd2751:BCD_Out <= 12'b000101101000;
		12'd2752:BCD_Out <= 12'b000101101000;
		12'd2753:BCD_Out <= 12'b000101101000;
		12'd2754:BCD_Out <= 12'b000101101000;
		12'd2755:BCD_Out <= 12'b000101101000;
		12'd2756:BCD_Out <= 12'b000101101000;
		12'd2757:BCD_Out <= 12'b000101101000;
		12'd2758:BCD_Out <= 12'b000101101000;
		12'd2759:BCD_Out <= 12'b000101101000;
		12'd2760:BCD_Out <= 12'b000101101000;
		12'd2761:BCD_Out <= 12'b000101101001;
		12'd2762:BCD_Out <= 12'b000101101001;
		12'd2763:BCD_Out <= 12'b000101101001;
		12'd2764:BCD_Out <= 12'b000101101001;
		12'd2765:BCD_Out <= 12'b000101101001;
		12'd2766:BCD_Out <= 12'b000101101001;
		12'd2767:BCD_Out <= 12'b000101101001;
		12'd2768:BCD_Out <= 12'b000101101001;
		12'd2769:BCD_Out <= 12'b000101101001;
		12'd2770:BCD_Out <= 12'b000101101001;
		12'd2771:BCD_Out <= 12'b000101101001;
		12'd2772:BCD_Out <= 12'b000101101001;
		12'd2773:BCD_Out <= 12'b000101101001;
		12'd2774:BCD_Out <= 12'b000101101001;
		12'd2775:BCD_Out <= 12'b000101101001;
		12'd2776:BCD_Out <= 12'b000101101001;
		12'd2777:BCD_Out <= 12'b000101110000;
		12'd2778:BCD_Out <= 12'b000101110000;
		12'd2779:BCD_Out <= 12'b000101110000;
		12'd2780:BCD_Out <= 12'b000101110000;
		12'd2781:BCD_Out <= 12'b000101110000;
		12'd2782:BCD_Out <= 12'b000101110000;
		12'd2783:BCD_Out <= 12'b000101110000;
		12'd2784:BCD_Out <= 12'b000101110000;
		12'd2785:BCD_Out <= 12'b000101110000;
		12'd2786:BCD_Out <= 12'b000101110000;
		12'd2787:BCD_Out <= 12'b000101110000;
		12'd2788:BCD_Out <= 12'b000101110000;
		12'd2789:BCD_Out <= 12'b000101110000;
		12'd2790:BCD_Out <= 12'b000101110000;
		12'd2791:BCD_Out <= 12'b000101110000;
		12'd2792:BCD_Out <= 12'b000101110000;
		12'd2793:BCD_Out <= 12'b000101110001;
		12'd2794:BCD_Out <= 12'b000101110001;
		12'd2795:BCD_Out <= 12'b000101110001;
		12'd2796:BCD_Out <= 12'b000101110001;
		12'd2797:BCD_Out <= 12'b000101110001;
		12'd2798:BCD_Out <= 12'b000101110001;
		12'd2799:BCD_Out <= 12'b000101110001;
		12'd2800:BCD_Out <= 12'b000101110001;
		12'd2801:BCD_Out <= 12'b000101110001;
		12'd2802:BCD_Out <= 12'b000101110001;
		12'd2803:BCD_Out <= 12'b000101110001;
		12'd2804:BCD_Out <= 12'b000101110001;
		12'd2805:BCD_Out <= 12'b000101110001;
		12'd2806:BCD_Out <= 12'b000101110001;
		12'd2807:BCD_Out <= 12'b000101110001;
		12'd2808:BCD_Out <= 12'b000101110001;
		12'd2809:BCD_Out <= 12'b000101110001;
		12'd2810:BCD_Out <= 12'b000101110010;
		12'd2811:BCD_Out <= 12'b000101110010;
		12'd2812:BCD_Out <= 12'b000101110010;
		12'd2813:BCD_Out <= 12'b000101110010;
		12'd2814:BCD_Out <= 12'b000101110010;
		12'd2815:BCD_Out <= 12'b000101110010;
		12'd2816:BCD_Out <= 12'b000101110010;
		12'd2817:BCD_Out <= 12'b000101110010;
		12'd2818:BCD_Out <= 12'b000101110010;
		12'd2819:BCD_Out <= 12'b000101110010;
		12'd2820:BCD_Out <= 12'b000101110010;
		12'd2821:BCD_Out <= 12'b000101110010;
		12'd2822:BCD_Out <= 12'b000101110010;
		12'd2823:BCD_Out <= 12'b000101110010;
		12'd2824:BCD_Out <= 12'b000101110010;
		12'd2825:BCD_Out <= 12'b000101110010;
		12'd2826:BCD_Out <= 12'b000101110011;
		12'd2827:BCD_Out <= 12'b000101110011;
		12'd2828:BCD_Out <= 12'b000101110011;
		12'd2829:BCD_Out <= 12'b000101110011;
		12'd2830:BCD_Out <= 12'b000101110011;
		12'd2831:BCD_Out <= 12'b000101110011;
		12'd2832:BCD_Out <= 12'b000101110011;
		12'd2833:BCD_Out <= 12'b000101110011;
		12'd2834:BCD_Out <= 12'b000101110011;
		12'd2835:BCD_Out <= 12'b000101110011;
		12'd2836:BCD_Out <= 12'b000101110011;
		12'd2837:BCD_Out <= 12'b000101110011;
		12'd2838:BCD_Out <= 12'b000101110011;
		12'd2839:BCD_Out <= 12'b000101110011;
		12'd2840:BCD_Out <= 12'b000101110011;
		12'd2841:BCD_Out <= 12'b000101110011;
		12'd2842:BCD_Out <= 12'b000101110100;
		12'd2843:BCD_Out <= 12'b000101110100;
		12'd2844:BCD_Out <= 12'b000101110100;
		12'd2845:BCD_Out <= 12'b000101110100;
		12'd2846:BCD_Out <= 12'b000101110100;
		12'd2847:BCD_Out <= 12'b000101110100;
		12'd2848:BCD_Out <= 12'b000101110100;
		12'd2849:BCD_Out <= 12'b000101110100;
		12'd2850:BCD_Out <= 12'b000101110100;
		12'd2851:BCD_Out <= 12'b000101110100;
		12'd2852:BCD_Out <= 12'b000101110100;
		12'd2853:BCD_Out <= 12'b000101110100;
		12'd2854:BCD_Out <= 12'b000101110100;
		12'd2855:BCD_Out <= 12'b000101110100;
		12'd2856:BCD_Out <= 12'b000101110100;
		12'd2857:BCD_Out <= 12'b000101110100;
		12'd2858:BCD_Out <= 12'b000101110100;
		12'd2859:BCD_Out <= 12'b000101110101;
		12'd2860:BCD_Out <= 12'b000101110101;
		12'd2861:BCD_Out <= 12'b000101110101;
		12'd2862:BCD_Out <= 12'b000101110101;
		12'd2863:BCD_Out <= 12'b000101110101;
		12'd2864:BCD_Out <= 12'b000101110101;
		12'd2865:BCD_Out <= 12'b000101110101;
		12'd2866:BCD_Out <= 12'b000101110101;
		12'd2867:BCD_Out <= 12'b000101110101;
		12'd2868:BCD_Out <= 12'b000101110101;
		12'd2869:BCD_Out <= 12'b000101110101;
		12'd2870:BCD_Out <= 12'b000101110101;
		12'd2871:BCD_Out <= 12'b000101110101;
		12'd2872:BCD_Out <= 12'b000101110101;
		12'd2873:BCD_Out <= 12'b000101110101;
		12'd2874:BCD_Out <= 12'b000101110101;
		12'd2875:BCD_Out <= 12'b000101110110;
		12'd2876:BCD_Out <= 12'b000101110110;
		12'd2877:BCD_Out <= 12'b000101110110;
		12'd2878:BCD_Out <= 12'b000101110110;
		12'd2879:BCD_Out <= 12'b000101110110;
		12'd2880:BCD_Out <= 12'b000101110110;
		12'd2881:BCD_Out <= 12'b000101110110;
		12'd2882:BCD_Out <= 12'b000101110110;
		12'd2883:BCD_Out <= 12'b000101110110;
		12'd2884:BCD_Out <= 12'b000101110110;
		12'd2885:BCD_Out <= 12'b000101110110;
		12'd2886:BCD_Out <= 12'b000101110110;
		12'd2887:BCD_Out <= 12'b000101110110;
		12'd2888:BCD_Out <= 12'b000101110110;
		12'd2889:BCD_Out <= 12'b000101110110;
		12'd2890:BCD_Out <= 12'b000101110110;
		12'd2891:BCD_Out <= 12'b000101110110;
		12'd2892:BCD_Out <= 12'b000101110111;
		12'd2893:BCD_Out <= 12'b000101110111;
		12'd2894:BCD_Out <= 12'b000101110111;
		12'd2895:BCD_Out <= 12'b000101110111;
		12'd2896:BCD_Out <= 12'b000101110111;
		12'd2897:BCD_Out <= 12'b000101110111;
		12'd2898:BCD_Out <= 12'b000101110111;
		12'd2899:BCD_Out <= 12'b000101110111;
		12'd2900:BCD_Out <= 12'b000101110111;
		12'd2901:BCD_Out <= 12'b000101110111;
		12'd2902:BCD_Out <= 12'b000101110111;
		12'd2903:BCD_Out <= 12'b000101110111;
		12'd2904:BCD_Out <= 12'b000101110111;
		12'd2905:BCD_Out <= 12'b000101110111;
		12'd2906:BCD_Out <= 12'b000101110111;
		12'd2907:BCD_Out <= 12'b000101110111;
		12'd2908:BCD_Out <= 12'b000101111000;
		12'd2909:BCD_Out <= 12'b000101111000;
		12'd2910:BCD_Out <= 12'b000101111000;
		12'd2911:BCD_Out <= 12'b000101111000;
		12'd2912:BCD_Out <= 12'b000101111000;
		12'd2913:BCD_Out <= 12'b000101111000;
		12'd2914:BCD_Out <= 12'b000101111000;
		12'd2915:BCD_Out <= 12'b000101111000;
		12'd2916:BCD_Out <= 12'b000101111000;
		12'd2917:BCD_Out <= 12'b000101111000;
		12'd2918:BCD_Out <= 12'b000101111000;
		12'd2919:BCD_Out <= 12'b000101111000;
		12'd2920:BCD_Out <= 12'b000101111000;
		12'd2921:BCD_Out <= 12'b000101111000;
		12'd2922:BCD_Out <= 12'b000101111000;
		12'd2923:BCD_Out <= 12'b000101111000;
		12'd2924:BCD_Out <= 12'b000101111001;
		12'd2925:BCD_Out <= 12'b000101111001;
		12'd2926:BCD_Out <= 12'b000101111001;
		12'd2927:BCD_Out <= 12'b000101111001;
		12'd2928:BCD_Out <= 12'b000101111001;
		12'd2929:BCD_Out <= 12'b000101111001;
		12'd2930:BCD_Out <= 12'b000101111001;
		12'd2931:BCD_Out <= 12'b000101111001;
		12'd2932:BCD_Out <= 12'b000101111001;
		12'd2933:BCD_Out <= 12'b000101111001;
		12'd2934:BCD_Out <= 12'b000101111001;
		12'd2935:BCD_Out <= 12'b000101111001;
		12'd2936:BCD_Out <= 12'b000101111001;
		12'd2937:BCD_Out <= 12'b000101111001;
		12'd2938:BCD_Out <= 12'b000101111001;
		12'd2939:BCD_Out <= 12'b000101111001;
		12'd2940:BCD_Out <= 12'b000101111001;
		12'd2941:BCD_Out <= 12'b000110000000;
		12'd2942:BCD_Out <= 12'b000110000000;
		12'd2943:BCD_Out <= 12'b000110000000;
		12'd2944:BCD_Out <= 12'b000110000000;
		12'd2945:BCD_Out <= 12'b000110000000;
		12'd2946:BCD_Out <= 12'b000110000000;
		12'd2947:BCD_Out <= 12'b000110000000;
		12'd2948:BCD_Out <= 12'b000110000000;
		12'd2949:BCD_Out <= 12'b000110000000;
		12'd2950:BCD_Out <= 12'b000110000000;
		12'd2951:BCD_Out <= 12'b000110000000;
		12'd2952:BCD_Out <= 12'b000110000000;
		12'd2953:BCD_Out <= 12'b000110000000;
		12'd2954:BCD_Out <= 12'b000110000000;
		12'd2955:BCD_Out <= 12'b000110000000;
		12'd2956:BCD_Out <= 12'b000110000000;
		12'd2957:BCD_Out <= 12'b000110000001;
		12'd2958:BCD_Out <= 12'b000110000001;
		12'd2959:BCD_Out <= 12'b000110000001;
		12'd2960:BCD_Out <= 12'b000110000001;
		12'd2961:BCD_Out <= 12'b000110000001;
		12'd2962:BCD_Out <= 12'b000110000001;
		12'd2963:BCD_Out <= 12'b000110000001;
		12'd2964:BCD_Out <= 12'b000110000001;
		12'd2965:BCD_Out <= 12'b000110000001;
		12'd2966:BCD_Out <= 12'b000110000001;
		12'd2967:BCD_Out <= 12'b000110000001;
		12'd2968:BCD_Out <= 12'b000110000001;
		12'd2969:BCD_Out <= 12'b000110000001;
		12'd2970:BCD_Out <= 12'b000110000001;
		12'd2971:BCD_Out <= 12'b000110000001;
		12'd2972:BCD_Out <= 12'b000110000001;
		12'd2973:BCD_Out <= 12'b000110000010;
		12'd2974:BCD_Out <= 12'b000110000010;
		12'd2975:BCD_Out <= 12'b000110000010;
		12'd2976:BCD_Out <= 12'b000110000010;
		12'd2977:BCD_Out <= 12'b000110000010;
		12'd2978:BCD_Out <= 12'b000110000010;
		12'd2979:BCD_Out <= 12'b000110000010;
		12'd2980:BCD_Out <= 12'b000110000010;
		12'd2981:BCD_Out <= 12'b000110000010;
		12'd2982:BCD_Out <= 12'b000110000010;
		12'd2983:BCD_Out <= 12'b000110000010;
		12'd2984:BCD_Out <= 12'b000110000010;
		12'd2985:BCD_Out <= 12'b000110000010;
		12'd2986:BCD_Out <= 12'b000110000010;
		12'd2987:BCD_Out <= 12'b000110000010;
		12'd2988:BCD_Out <= 12'b000110000010;
		12'd2989:BCD_Out <= 12'b000110000010;
		12'd2990:BCD_Out <= 12'b000110000011;
		12'd2991:BCD_Out <= 12'b000110000011;
		12'd2992:BCD_Out <= 12'b000110000011;
		12'd2993:BCD_Out <= 12'b000110000011;
		12'd2994:BCD_Out <= 12'b000110000011;
		12'd2995:BCD_Out <= 12'b000110000011;
		12'd2996:BCD_Out <= 12'b000110000011;
		12'd2997:BCD_Out <= 12'b000110000011;
		12'd2998:BCD_Out <= 12'b000110000011;
		12'd2999:BCD_Out <= 12'b000110000011;
		12'd3000:BCD_Out <= 12'b000110000011;
		12'd3001:BCD_Out <= 12'b000110000011;
		12'd3002:BCD_Out <= 12'b000110000011;
		12'd3003:BCD_Out <= 12'b000110000011;
		12'd3004:BCD_Out <= 12'b000110000011;
		12'd3005:BCD_Out <= 12'b000110000011;
		12'd3006:BCD_Out <= 12'b000110000100;
		12'd3007:BCD_Out <= 12'b000110000100;
		12'd3008:BCD_Out <= 12'b000110000100;
		12'd3009:BCD_Out <= 12'b000110000100;
		12'd3010:BCD_Out <= 12'b000110000100;
		12'd3011:BCD_Out <= 12'b000110000100;
		12'd3012:BCD_Out <= 12'b000110000100;
		12'd3013:BCD_Out <= 12'b000110000100;
		12'd3014:BCD_Out <= 12'b000110000100;
		12'd3015:BCD_Out <= 12'b000110000100;
		12'd3016:BCD_Out <= 12'b000110000100;
		12'd3017:BCD_Out <= 12'b000110000100;
		12'd3018:BCD_Out <= 12'b000110000100;
		12'd3019:BCD_Out <= 12'b000110000100;
		12'd3020:BCD_Out <= 12'b000110000100;
		12'd3021:BCD_Out <= 12'b000110000100;
		12'd3022:BCD_Out <= 12'b000110000100;
		12'd3023:BCD_Out <= 12'b000110000101;
		12'd3024:BCD_Out <= 12'b000110000101;
		12'd3025:BCD_Out <= 12'b000110000101;
		12'd3026:BCD_Out <= 12'b000110000101;
		12'd3027:BCD_Out <= 12'b000110000101;
		12'd3028:BCD_Out <= 12'b000110000101;
		12'd3029:BCD_Out <= 12'b000110000101;
		12'd3030:BCD_Out <= 12'b000110000101;
		12'd3031:BCD_Out <= 12'b000110000101;
		12'd3032:BCD_Out <= 12'b000110000101;
		12'd3033:BCD_Out <= 12'b000110000101;
		12'd3034:BCD_Out <= 12'b000110000101;
		12'd3035:BCD_Out <= 12'b000110000101;
		12'd3036:BCD_Out <= 12'b000110000101;
		12'd3037:BCD_Out <= 12'b000110000101;
		12'd3038:BCD_Out <= 12'b000110000101;
		12'd3039:BCD_Out <= 12'b000110000110;
		12'd3040:BCD_Out <= 12'b000110000110;
		12'd3041:BCD_Out <= 12'b000110000110;
		12'd3042:BCD_Out <= 12'b000110000110;
		12'd3043:BCD_Out <= 12'b000110000110;
		12'd3044:BCD_Out <= 12'b000110000110;
		12'd3045:BCD_Out <= 12'b000110000110;
		12'd3046:BCD_Out <= 12'b000110000110;
		12'd3047:BCD_Out <= 12'b000110000110;
		12'd3048:BCD_Out <= 12'b000110000110;
		12'd3049:BCD_Out <= 12'b000110000110;
		12'd3050:BCD_Out <= 12'b000110000110;
		12'd3051:BCD_Out <= 12'b000110000110;
		12'd3052:BCD_Out <= 12'b000110000110;
		12'd3053:BCD_Out <= 12'b000110000110;
		12'd3054:BCD_Out <= 12'b000110000110;
		12'd3055:BCD_Out <= 12'b000110000111;
		12'd3056:BCD_Out <= 12'b000110000111;
		12'd3057:BCD_Out <= 12'b000110000111;
		12'd3058:BCD_Out <= 12'b000110000111;
		12'd3059:BCD_Out <= 12'b000110000111;
		12'd3060:BCD_Out <= 12'b000110000111;
		12'd3061:BCD_Out <= 12'b000110000111;
		12'd3062:BCD_Out <= 12'b000110000111;
		12'd3063:BCD_Out <= 12'b000110000111;
		12'd3064:BCD_Out <= 12'b000110000111;
		12'd3065:BCD_Out <= 12'b000110000111;
		12'd3066:BCD_Out <= 12'b000110000111;
		12'd3067:BCD_Out <= 12'b000110000111;
		12'd3068:BCD_Out <= 12'b000110000111;
		12'd3069:BCD_Out <= 12'b000110000111;
		12'd3070:BCD_Out <= 12'b000110000111;
		12'd3071:BCD_Out <= 12'b000110000111;
		12'd3072:BCD_Out <= 12'b000110001000;
		12'd3073:BCD_Out <= 12'b000110001000;
		12'd3074:BCD_Out <= 12'b000110001000;
		12'd3075:BCD_Out <= 12'b000110001000;
		12'd3076:BCD_Out <= 12'b000110001000;
		12'd3077:BCD_Out <= 12'b000110001000;
		12'd3078:BCD_Out <= 12'b000110001000;
		12'd3079:BCD_Out <= 12'b000110001000;
		12'd3080:BCD_Out <= 12'b000110001000;
		12'd3081:BCD_Out <= 12'b000110001000;
		12'd3082:BCD_Out <= 12'b000110001000;
		12'd3083:BCD_Out <= 12'b000110001000;
		12'd3084:BCD_Out <= 12'b000110001000;
		12'd3085:BCD_Out <= 12'b000110001000;
		12'd3086:BCD_Out <= 12'b000110001000;
		12'd3087:BCD_Out <= 12'b000110001000;
		12'd3088:BCD_Out <= 12'b000110001001;
		12'd3089:BCD_Out <= 12'b000110001001;
		12'd3090:BCD_Out <= 12'b000110001001;
		12'd3091:BCD_Out <= 12'b000110001001;
		12'd3092:BCD_Out <= 12'b000110001001;
		12'd3093:BCD_Out <= 12'b000110001001;
		12'd3094:BCD_Out <= 12'b000110001001;
		12'd3095:BCD_Out <= 12'b000110001001;
		12'd3096:BCD_Out <= 12'b000110001001;
		12'd3097:BCD_Out <= 12'b000110001001;
		12'd3098:BCD_Out <= 12'b000110001001;
		12'd3099:BCD_Out <= 12'b000110001001;
		12'd3100:BCD_Out <= 12'b000110001001;
		12'd3101:BCD_Out <= 12'b000110001001;
		12'd3102:BCD_Out <= 12'b000110001001;
		12'd3103:BCD_Out <= 12'b000110001001;
		12'd3104:BCD_Out <= 12'b000110001001;
		12'd3105:BCD_Out <= 12'b000110010000;
		12'd3106:BCD_Out <= 12'b000110010000;
		12'd3107:BCD_Out <= 12'b000110010000;
		12'd3108:BCD_Out <= 12'b000110010000;
		12'd3109:BCD_Out <= 12'b000110010000;
		12'd3110:BCD_Out <= 12'b000110010000;
		12'd3111:BCD_Out <= 12'b000110010000;
		12'd3112:BCD_Out <= 12'b000110010000;
		12'd3113:BCD_Out <= 12'b000110010000;
		12'd3114:BCD_Out <= 12'b000110010000;
		12'd3115:BCD_Out <= 12'b000110010000;
		12'd3116:BCD_Out <= 12'b000110010000;
		12'd3117:BCD_Out <= 12'b000110010000;
		12'd3118:BCD_Out <= 12'b000110010000;
		12'd3119:BCD_Out <= 12'b000110010000;
		12'd3120:BCD_Out <= 12'b000110010000;
		12'd3121:BCD_Out <= 12'b000110010001;
		12'd3122:BCD_Out <= 12'b000110010001;
		12'd3123:BCD_Out <= 12'b000110010001;
		12'd3124:BCD_Out <= 12'b000110010001;
		12'd3125:BCD_Out <= 12'b000110010001;
		12'd3126:BCD_Out <= 12'b000110010001;
		12'd3127:BCD_Out <= 12'b000110010001;
		12'd3128:BCD_Out <= 12'b000110010001;
		12'd3129:BCD_Out <= 12'b000110010001;
		12'd3130:BCD_Out <= 12'b000110010001;
		12'd3131:BCD_Out <= 12'b000110010001;
		12'd3132:BCD_Out <= 12'b000110010001;
		12'd3133:BCD_Out <= 12'b000110010001;
		12'd3134:BCD_Out <= 12'b000110010001;
		12'd3135:BCD_Out <= 12'b000110010001;
		12'd3136:BCD_Out <= 12'b000110010001;
		12'd3137:BCD_Out <= 12'b000110010010;
		12'd3138:BCD_Out <= 12'b000110010010;
		12'd3139:BCD_Out <= 12'b000110010010;
		12'd3140:BCD_Out <= 12'b000110010010;
		12'd3141:BCD_Out <= 12'b000110010010;
		12'd3142:BCD_Out <= 12'b000110010010;
		12'd3143:BCD_Out <= 12'b000110010010;
		12'd3144:BCD_Out <= 12'b000110010010;
		12'd3145:BCD_Out <= 12'b000110010010;
		12'd3146:BCD_Out <= 12'b000110010010;
		12'd3147:BCD_Out <= 12'b000110010010;
		12'd3148:BCD_Out <= 12'b000110010010;
		12'd3149:BCD_Out <= 12'b000110010010;
		12'd3150:BCD_Out <= 12'b000110010010;
		12'd3151:BCD_Out <= 12'b000110010010;
		12'd3152:BCD_Out <= 12'b000110010010;
		12'd3153:BCD_Out <= 12'b000110010010;
		12'd3154:BCD_Out <= 12'b000110010011;
		12'd3155:BCD_Out <= 12'b000110010011;
		12'd3156:BCD_Out <= 12'b000110010011;
		12'd3157:BCD_Out <= 12'b000110010011;
		12'd3158:BCD_Out <= 12'b000110010011;
		12'd3159:BCD_Out <= 12'b000110010011;
		12'd3160:BCD_Out <= 12'b000110010011;
		12'd3161:BCD_Out <= 12'b000110010011;
		12'd3162:BCD_Out <= 12'b000110010011;
		12'd3163:BCD_Out <= 12'b000110010011;
		12'd3164:BCD_Out <= 12'b000110010011;
		12'd3165:BCD_Out <= 12'b000110010011;
		12'd3166:BCD_Out <= 12'b000110010011;
		12'd3167:BCD_Out <= 12'b000110010011;
		12'd3168:BCD_Out <= 12'b000110010011;
		12'd3169:BCD_Out <= 12'b000110010011;
		12'd3170:BCD_Out <= 12'b000110010100;
		12'd3171:BCD_Out <= 12'b000110010100;
		12'd3172:BCD_Out <= 12'b000110010100;
		12'd3173:BCD_Out <= 12'b000110010100;
		12'd3174:BCD_Out <= 12'b000110010100;
		12'd3175:BCD_Out <= 12'b000110010100;
		12'd3176:BCD_Out <= 12'b000110010100;
		12'd3177:BCD_Out <= 12'b000110010100;
		12'd3178:BCD_Out <= 12'b000110010100;
		12'd3179:BCD_Out <= 12'b000110010100;
		12'd3180:BCD_Out <= 12'b000110010100;
		12'd3181:BCD_Out <= 12'b000110010100;
		12'd3182:BCD_Out <= 12'b000110010100;
		12'd3183:BCD_Out <= 12'b000110010100;
		12'd3184:BCD_Out <= 12'b000110010100;
		12'd3185:BCD_Out <= 12'b000110010100;
		12'd3186:BCD_Out <= 12'b000110010101;
		12'd3187:BCD_Out <= 12'b000110010101;
		12'd3188:BCD_Out <= 12'b000110010101;
		12'd3189:BCD_Out <= 12'b000110010101;
		12'd3190:BCD_Out <= 12'b000110010101;
		12'd3191:BCD_Out <= 12'b000110010101;
		12'd3192:BCD_Out <= 12'b000110010101;
		12'd3193:BCD_Out <= 12'b000110010101;
		12'd3194:BCD_Out <= 12'b000110010101;
		12'd3195:BCD_Out <= 12'b000110010101;
		12'd3196:BCD_Out <= 12'b000110010101;
		12'd3197:BCD_Out <= 12'b000110010101;
		12'd3198:BCD_Out <= 12'b000110010101;
		12'd3199:BCD_Out <= 12'b000110010101;
		12'd3200:BCD_Out <= 12'b000110010101;
		12'd3201:BCD_Out <= 12'b000110010101;
		12'd3202:BCD_Out <= 12'b000110010101;
		12'd3203:BCD_Out <= 12'b000110010110;
		12'd3204:BCD_Out <= 12'b000110010110;
		12'd3205:BCD_Out <= 12'b000110010110;
		12'd3206:BCD_Out <= 12'b000110010110;
		12'd3207:BCD_Out <= 12'b000110010110;
		12'd3208:BCD_Out <= 12'b000110010110;
		12'd3209:BCD_Out <= 12'b000110010110;
		12'd3210:BCD_Out <= 12'b000110010110;
		12'd3211:BCD_Out <= 12'b000110010110;
		12'd3212:BCD_Out <= 12'b000110010110;
		12'd3213:BCD_Out <= 12'b000110010110;
		12'd3214:BCD_Out <= 12'b000110010110;
		12'd3215:BCD_Out <= 12'b000110010110;
		12'd3216:BCD_Out <= 12'b000110010110;
		12'd3217:BCD_Out <= 12'b000110010110;
		12'd3218:BCD_Out <= 12'b000110010110;
		12'd3219:BCD_Out <= 12'b000110010111;
		12'd3220:BCD_Out <= 12'b000110010111;
		12'd3221:BCD_Out <= 12'b000110010111;
		12'd3222:BCD_Out <= 12'b000110010111;
		12'd3223:BCD_Out <= 12'b000110010111;
		12'd3224:BCD_Out <= 12'b000110010111;
		12'd3225:BCD_Out <= 12'b000110010111;
		12'd3226:BCD_Out <= 12'b000110010111;
		12'd3227:BCD_Out <= 12'b000110010111;
		12'd3228:BCD_Out <= 12'b000110010111;
		12'd3229:BCD_Out <= 12'b000110010111;
		12'd3230:BCD_Out <= 12'b000110010111;
		12'd3231:BCD_Out <= 12'b000110010111;
		12'd3232:BCD_Out <= 12'b000110010111;
		12'd3233:BCD_Out <= 12'b000110010111;
		12'd3234:BCD_Out <= 12'b000110010111;
		12'd3235:BCD_Out <= 12'b000110010111;
		12'd3236:BCD_Out <= 12'b000110011000;
		12'd3237:BCD_Out <= 12'b000110011000;
		12'd3238:BCD_Out <= 12'b000110011000;
		12'd3239:BCD_Out <= 12'b000110011000;
		12'd3240:BCD_Out <= 12'b000110011000;
		12'd3241:BCD_Out <= 12'b000110011000;
		12'd3242:BCD_Out <= 12'b000110011000;
		12'd3243:BCD_Out <= 12'b000110011000;
		12'd3244:BCD_Out <= 12'b000110011000;
		12'd3245:BCD_Out <= 12'b000110011000;
		12'd3246:BCD_Out <= 12'b000110011000;
		12'd3247:BCD_Out <= 12'b000110011000;
		12'd3248:BCD_Out <= 12'b000110011000;
		12'd3249:BCD_Out <= 12'b000110011000;
		12'd3250:BCD_Out <= 12'b000110011000;
		12'd3251:BCD_Out <= 12'b000110011000;
		12'd3252:BCD_Out <= 12'b000110011001;
		12'd3253:BCD_Out <= 12'b000110011001;
		12'd3254:BCD_Out <= 12'b000110011001;
		12'd3255:BCD_Out <= 12'b000110011001;
		12'd3256:BCD_Out <= 12'b000110011001;
		12'd3257:BCD_Out <= 12'b000110011001;
		12'd3258:BCD_Out <= 12'b000110011001;
		12'd3259:BCD_Out <= 12'b000110011001;
		12'd3260:BCD_Out <= 12'b000110011001;
		12'd3261:BCD_Out <= 12'b000110011001;
		12'd3262:BCD_Out <= 12'b000110011001;
		12'd3263:BCD_Out <= 12'b000110011001;
		12'd3264:BCD_Out <= 12'b000110011001;
		12'd3265:BCD_Out <= 12'b000110011001;
		12'd3266:BCD_Out <= 12'b000110011001;
		12'd3267:BCD_Out <= 12'b000110011001;
		12'd3268:BCD_Out <= 12'b001000000000;
		12'd3269:BCD_Out <= 12'b001000000000;
		12'd3270:BCD_Out <= 12'b001000000000;
		12'd3271:BCD_Out <= 12'b001000000000;
		12'd3272:BCD_Out <= 12'b001000000000;
		12'd3273:BCD_Out <= 12'b001000000000;
		12'd3274:BCD_Out <= 12'b001000000000;
		12'd3275:BCD_Out <= 12'b001000000000;
		12'd3276:BCD_Out <= 12'b001000000000;
		12'd3277:BCD_Out <= 12'b001000000000;
		12'd3278:BCD_Out <= 12'b001000000000;
		12'd3279:BCD_Out <= 12'b001000000000;
		12'd3280:BCD_Out <= 12'b001000000000;
		12'd3281:BCD_Out <= 12'b001000000000;
		12'd3282:BCD_Out <= 12'b001000000000;
		12'd3283:BCD_Out <= 12'b001000000000;
		12'd3284:BCD_Out <= 12'b001000000000;
		12'd3285:BCD_Out <= 12'b001000000001;
		12'd3286:BCD_Out <= 12'b001000000001;
		12'd3287:BCD_Out <= 12'b001000000001;
		12'd3288:BCD_Out <= 12'b001000000001;
		12'd3289:BCD_Out <= 12'b001000000001;
		12'd3290:BCD_Out <= 12'b001000000001;
		12'd3291:BCD_Out <= 12'b001000000001;
		12'd3292:BCD_Out <= 12'b001000000001;
		12'd3293:BCD_Out <= 12'b001000000001;
		12'd3294:BCD_Out <= 12'b001000000001;
		12'd3295:BCD_Out <= 12'b001000000001;
		12'd3296:BCD_Out <= 12'b001000000001;
		12'd3297:BCD_Out <= 12'b001000000001;
		12'd3298:BCD_Out <= 12'b001000000001;
		12'd3299:BCD_Out <= 12'b001000000001;
		12'd3300:BCD_Out <= 12'b001000000001;
		12'd3301:BCD_Out <= 12'b001000000010;
		12'd3302:BCD_Out <= 12'b001000000010;
		12'd3303:BCD_Out <= 12'b001000000010;
		12'd3304:BCD_Out <= 12'b001000000010;
		12'd3305:BCD_Out <= 12'b001000000010;
		12'd3306:BCD_Out <= 12'b001000000010;
		12'd3307:BCD_Out <= 12'b001000000010;
		12'd3308:BCD_Out <= 12'b001000000010;
		12'd3309:BCD_Out <= 12'b001000000010;
		12'd3310:BCD_Out <= 12'b001000000010;
		12'd3311:BCD_Out <= 12'b001000000010;
		12'd3312:BCD_Out <= 12'b001000000010;
		12'd3313:BCD_Out <= 12'b001000000010;
		12'd3314:BCD_Out <= 12'b001000000010;
		12'd3315:BCD_Out <= 12'b001000000010;
		12'd3316:BCD_Out <= 12'b001000000010;
		12'd3317:BCD_Out <= 12'b001000000011;
		12'd3318:BCD_Out <= 12'b001000000011;
		12'd3319:BCD_Out <= 12'b001000000011;
		12'd3320:BCD_Out <= 12'b001000000011;
		12'd3321:BCD_Out <= 12'b001000000011;
		12'd3322:BCD_Out <= 12'b001000000011;
		12'd3323:BCD_Out <= 12'b001000000011;
		12'd3324:BCD_Out <= 12'b001000000011;
		12'd3325:BCD_Out <= 12'b001000000011;
		12'd3326:BCD_Out <= 12'b001000000011;
		12'd3327:BCD_Out <= 12'b001000000011;
		12'd3328:BCD_Out <= 12'b001000000011;
		12'd3329:BCD_Out <= 12'b001000000011;
		12'd3330:BCD_Out <= 12'b001000000011;
		12'd3331:BCD_Out <= 12'b001000000011;
		12'd3332:BCD_Out <= 12'b001000000011;
		12'd3333:BCD_Out <= 12'b001000000011;
		12'd3334:BCD_Out <= 12'b001000000100;
		12'd3335:BCD_Out <= 12'b001000000100;
		12'd3336:BCD_Out <= 12'b001000000100;
		12'd3337:BCD_Out <= 12'b001000000100;
		12'd3338:BCD_Out <= 12'b001000000100;
		12'd3339:BCD_Out <= 12'b001000000100;
		12'd3340:BCD_Out <= 12'b001000000100;
		12'd3341:BCD_Out <= 12'b001000000100;
		12'd3342:BCD_Out <= 12'b001000000100;
		12'd3343:BCD_Out <= 12'b001000000100;
		12'd3344:BCD_Out <= 12'b001000000100;
		12'd3345:BCD_Out <= 12'b001000000100;
		12'd3346:BCD_Out <= 12'b001000000100;
		12'd3347:BCD_Out <= 12'b001000000100;
		12'd3348:BCD_Out <= 12'b001000000100;
		12'd3349:BCD_Out <= 12'b001000000100;
		12'd3350:BCD_Out <= 12'b001000000101;
		12'd3351:BCD_Out <= 12'b001000000101;
		12'd3352:BCD_Out <= 12'b001000000101;
		12'd3353:BCD_Out <= 12'b001000000101;
		12'd3354:BCD_Out <= 12'b001000000101;
		12'd3355:BCD_Out <= 12'b001000000101;
		12'd3356:BCD_Out <= 12'b001000000101;
		12'd3357:BCD_Out <= 12'b001000000101;
		12'd3358:BCD_Out <= 12'b001000000101;
		12'd3359:BCD_Out <= 12'b001000000101;
		12'd3360:BCD_Out <= 12'b001000000101;
		12'd3361:BCD_Out <= 12'b001000000101;
		12'd3362:BCD_Out <= 12'b001000000101;
		12'd3363:BCD_Out <= 12'b001000000101;
		12'd3364:BCD_Out <= 12'b001000000101;
		12'd3365:BCD_Out <= 12'b001000000101;
		12'd3366:BCD_Out <= 12'b001000000101;
		12'd3367:BCD_Out <= 12'b001000000110;
		12'd3368:BCD_Out <= 12'b001000000110;
		12'd3369:BCD_Out <= 12'b001000000110;
		12'd3370:BCD_Out <= 12'b001000000110;
		12'd3371:BCD_Out <= 12'b001000000110;
		12'd3372:BCD_Out <= 12'b001000000110;
		12'd3373:BCD_Out <= 12'b001000000110;
		12'd3374:BCD_Out <= 12'b001000000110;
		12'd3375:BCD_Out <= 12'b001000000110;
		12'd3376:BCD_Out <= 12'b001000000110;
		12'd3377:BCD_Out <= 12'b001000000110;
		12'd3378:BCD_Out <= 12'b001000000110;
		12'd3379:BCD_Out <= 12'b001000000110;
		12'd3380:BCD_Out <= 12'b001000000110;
		12'd3381:BCD_Out <= 12'b001000000110;
		12'd3382:BCD_Out <= 12'b001000000110;
		12'd3383:BCD_Out <= 12'b001000000111;
		12'd3384:BCD_Out <= 12'b001000000111;
		12'd3385:BCD_Out <= 12'b001000000111;
		12'd3386:BCD_Out <= 12'b001000000111;
		12'd3387:BCD_Out <= 12'b001000000111;
		12'd3388:BCD_Out <= 12'b001000000111;
		12'd3389:BCD_Out <= 12'b001000000111;
		12'd3390:BCD_Out <= 12'b001000000111;
		12'd3391:BCD_Out <= 12'b001000000111;
		12'd3392:BCD_Out <= 12'b001000000111;
		12'd3393:BCD_Out <= 12'b001000000111;
		12'd3394:BCD_Out <= 12'b001000000111;
		12'd3395:BCD_Out <= 12'b001000000111;
		12'd3396:BCD_Out <= 12'b001000000111;
		12'd3397:BCD_Out <= 12'b001000000111;
		12'd3398:BCD_Out <= 12'b001000000111;
		12'd3399:BCD_Out <= 12'b001000001000;
		12'd3400:BCD_Out <= 12'b001000001000;
		12'd3401:BCD_Out <= 12'b001000001000;
		12'd3402:BCD_Out <= 12'b001000001000;
		12'd3403:BCD_Out <= 12'b001000001000;
		12'd3404:BCD_Out <= 12'b001000001000;
		12'd3405:BCD_Out <= 12'b001000001000;
		12'd3406:BCD_Out <= 12'b001000001000;
		12'd3407:BCD_Out <= 12'b001000001000;
		12'd3408:BCD_Out <= 12'b001000001000;
		12'd3409:BCD_Out <= 12'b001000001000;
		12'd3410:BCD_Out <= 12'b001000001000;
		12'd3411:BCD_Out <= 12'b001000001000;
		12'd3412:BCD_Out <= 12'b001000001000;
		12'd3413:BCD_Out <= 12'b001000001000;
		12'd3414:BCD_Out <= 12'b001000001000;
		12'd3415:BCD_Out <= 12'b001000001000;
		12'd3416:BCD_Out <= 12'b001000001001;
		12'd3417:BCD_Out <= 12'b001000001001;
		12'd3418:BCD_Out <= 12'b001000001001;
		12'd3419:BCD_Out <= 12'b001000001001;
		12'd3420:BCD_Out <= 12'b001000001001;
		12'd3421:BCD_Out <= 12'b001000001001;
		12'd3422:BCD_Out <= 12'b001000001001;
		12'd3423:BCD_Out <= 12'b001000001001;
		12'd3424:BCD_Out <= 12'b001000001001;
		12'd3425:BCD_Out <= 12'b001000001001;
		12'd3426:BCD_Out <= 12'b001000001001;
		12'd3427:BCD_Out <= 12'b001000001001;
		12'd3428:BCD_Out <= 12'b001000001001;
		12'd3429:BCD_Out <= 12'b001000001001;
		12'd3430:BCD_Out <= 12'b001000001001;
		12'd3431:BCD_Out <= 12'b001000001001;
		12'd3432:BCD_Out <= 12'b001000010000;
		12'd3433:BCD_Out <= 12'b001000010000;
		12'd3434:BCD_Out <= 12'b001000010000;
		12'd3435:BCD_Out <= 12'b001000010000;
		12'd3436:BCD_Out <= 12'b001000010000;
		12'd3437:BCD_Out <= 12'b001000010000;
		12'd3438:BCD_Out <= 12'b001000010000;
		12'd3439:BCD_Out <= 12'b001000010000;
		12'd3440:BCD_Out <= 12'b001000010000;
		12'd3441:BCD_Out <= 12'b001000010000;
		12'd3442:BCD_Out <= 12'b001000010000;
		12'd3443:BCD_Out <= 12'b001000010000;
		12'd3444:BCD_Out <= 12'b001000010000;
		12'd3445:BCD_Out <= 12'b001000010000;
		12'd3446:BCD_Out <= 12'b001000010000;
		12'd3447:BCD_Out <= 12'b001000010000;
		12'd3448:BCD_Out <= 12'b001000010001;
		12'd3449:BCD_Out <= 12'b001000010001;
		12'd3450:BCD_Out <= 12'b001000010001;
		12'd3451:BCD_Out <= 12'b001000010001;
		12'd3452:BCD_Out <= 12'b001000010001;
		12'd3453:BCD_Out <= 12'b001000010001;
		12'd3454:BCD_Out <= 12'b001000010001;
		12'd3455:BCD_Out <= 12'b001000010001;
		12'd3456:BCD_Out <= 12'b001000010001;
		12'd3457:BCD_Out <= 12'b001000010001;
		12'd3458:BCD_Out <= 12'b001000010001;
		12'd3459:BCD_Out <= 12'b001000010001;
		12'd3460:BCD_Out <= 12'b001000010001;
		12'd3461:BCD_Out <= 12'b001000010001;
		12'd3462:BCD_Out <= 12'b001000010001;
		12'd3463:BCD_Out <= 12'b001000010001;
		12'd3464:BCD_Out <= 12'b001000010001;
		12'd3465:BCD_Out <= 12'b001000010010;
		12'd3466:BCD_Out <= 12'b001000010010;
		12'd3467:BCD_Out <= 12'b001000010010;
		12'd3468:BCD_Out <= 12'b001000010010;
		12'd3469:BCD_Out <= 12'b001000010010;
		12'd3470:BCD_Out <= 12'b001000010010;
		12'd3471:BCD_Out <= 12'b001000010010;
		12'd3472:BCD_Out <= 12'b001000010010;
		12'd3473:BCD_Out <= 12'b001000010010;
		12'd3474:BCD_Out <= 12'b001000010010;
		12'd3475:BCD_Out <= 12'b001000010010;
		12'd3476:BCD_Out <= 12'b001000010010;
		12'd3477:BCD_Out <= 12'b001000010010;
		12'd3478:BCD_Out <= 12'b001000010010;
		12'd3479:BCD_Out <= 12'b001000010010;
		12'd3480:BCD_Out <= 12'b001000010010;
		12'd3481:BCD_Out <= 12'b001000010011;
		12'd3482:BCD_Out <= 12'b001000010011;
		12'd3483:BCD_Out <= 12'b001000010011;
		12'd3484:BCD_Out <= 12'b001000010011;
		12'd3485:BCD_Out <= 12'b001000010011;
		12'd3486:BCD_Out <= 12'b001000010011;
		12'd3487:BCD_Out <= 12'b001000010011;
		12'd3488:BCD_Out <= 12'b001000010011;
		12'd3489:BCD_Out <= 12'b001000010011;
		12'd3490:BCD_Out <= 12'b001000010011;
		12'd3491:BCD_Out <= 12'b001000010011;
		12'd3492:BCD_Out <= 12'b001000010011;
		12'd3493:BCD_Out <= 12'b001000010011;
		12'd3494:BCD_Out <= 12'b001000010011;
		12'd3495:BCD_Out <= 12'b001000010011;
		12'd3496:BCD_Out <= 12'b001000010011;
		12'd3497:BCD_Out <= 12'b001000010011;
		12'd3498:BCD_Out <= 12'b001000010100;
		12'd3499:BCD_Out <= 12'b001000010100;
		12'd3500:BCD_Out <= 12'b001000010100;
		12'd3501:BCD_Out <= 12'b001000010100;
		12'd3502:BCD_Out <= 12'b001000010100;
		12'd3503:BCD_Out <= 12'b001000010100;
		12'd3504:BCD_Out <= 12'b001000010100;
		12'd3505:BCD_Out <= 12'b001000010100;
		12'd3506:BCD_Out <= 12'b001000010100;
		12'd3507:BCD_Out <= 12'b001000010100;
		12'd3508:BCD_Out <= 12'b001000010100;
		12'd3509:BCD_Out <= 12'b001000010100;
		12'd3510:BCD_Out <= 12'b001000010100;
		12'd3511:BCD_Out <= 12'b001000010100;
		12'd3512:BCD_Out <= 12'b001000010100;
		12'd3513:BCD_Out <= 12'b001000010100;
		12'd3514:BCD_Out <= 12'b001000010101;
		12'd3515:BCD_Out <= 12'b001000010101;
		12'd3516:BCD_Out <= 12'b001000010101;
		12'd3517:BCD_Out <= 12'b001000010101;
		12'd3518:BCD_Out <= 12'b001000010101;
		12'd3519:BCD_Out <= 12'b001000010101;
		12'd3520:BCD_Out <= 12'b001000010101;
		12'd3521:BCD_Out <= 12'b001000010101;
		12'd3522:BCD_Out <= 12'b001000010101;
		12'd3523:BCD_Out <= 12'b001000010101;
		12'd3524:BCD_Out <= 12'b001000010101;
		12'd3525:BCD_Out <= 12'b001000010101;
		12'd3526:BCD_Out <= 12'b001000010101;
		12'd3527:BCD_Out <= 12'b001000010101;
		12'd3528:BCD_Out <= 12'b001000010101;
		12'd3529:BCD_Out <= 12'b001000010101;
		12'd3530:BCD_Out <= 12'b001000010110;
		12'd3531:BCD_Out <= 12'b001000010110;
		12'd3532:BCD_Out <= 12'b001000010110;
		12'd3533:BCD_Out <= 12'b001000010110;
		12'd3534:BCD_Out <= 12'b001000010110;
		12'd3535:BCD_Out <= 12'b001000010110;
		12'd3536:BCD_Out <= 12'b001000010110;
		12'd3537:BCD_Out <= 12'b001000010110;
		12'd3538:BCD_Out <= 12'b001000010110;
		12'd3539:BCD_Out <= 12'b001000010110;
		12'd3540:BCD_Out <= 12'b001000010110;
		12'd3541:BCD_Out <= 12'b001000010110;
		12'd3542:BCD_Out <= 12'b001000010110;
		12'd3543:BCD_Out <= 12'b001000010110;
		12'd3544:BCD_Out <= 12'b001000010110;
		12'd3545:BCD_Out <= 12'b001000010110;
		12'd3546:BCD_Out <= 12'b001000010110;
		12'd3547:BCD_Out <= 12'b001000010111;
		12'd3548:BCD_Out <= 12'b001000010111;
		12'd3549:BCD_Out <= 12'b001000010111;
		12'd3550:BCD_Out <= 12'b001000010111;
		12'd3551:BCD_Out <= 12'b001000010111;
		12'd3552:BCD_Out <= 12'b001000010111;
		12'd3553:BCD_Out <= 12'b001000010111;
		12'd3554:BCD_Out <= 12'b001000010111;
		12'd3555:BCD_Out <= 12'b001000010111;
		12'd3556:BCD_Out <= 12'b001000010111;
		12'd3557:BCD_Out <= 12'b001000010111;
		12'd3558:BCD_Out <= 12'b001000010111;
		12'd3559:BCD_Out <= 12'b001000010111;
		12'd3560:BCD_Out <= 12'b001000010111;
		12'd3561:BCD_Out <= 12'b001000010111;
		12'd3562:BCD_Out <= 12'b001000010111;
		12'd3563:BCD_Out <= 12'b001000011000;
		12'd3564:BCD_Out <= 12'b001000011000;
		12'd3565:BCD_Out <= 12'b001000011000;
		12'd3566:BCD_Out <= 12'b001000011000;
		12'd3567:BCD_Out <= 12'b001000011000;
		12'd3568:BCD_Out <= 12'b001000011000;
		12'd3569:BCD_Out <= 12'b001000011000;
		12'd3570:BCD_Out <= 12'b001000011000;
		12'd3571:BCD_Out <= 12'b001000011000;
		12'd3572:BCD_Out <= 12'b001000011000;
		12'd3573:BCD_Out <= 12'b001000011000;
		12'd3574:BCD_Out <= 12'b001000011000;
		12'd3575:BCD_Out <= 12'b001000011000;
		12'd3576:BCD_Out <= 12'b001000011000;
		12'd3577:BCD_Out <= 12'b001000011000;
		12'd3578:BCD_Out <= 12'b001000011000;
		12'd3579:BCD_Out <= 12'b001000011000;
		12'd3580:BCD_Out <= 12'b001000011001;
		12'd3581:BCD_Out <= 12'b001000011001;
		12'd3582:BCD_Out <= 12'b001000011001;
		12'd3583:BCD_Out <= 12'b001000011001;
		12'd3584:BCD_Out <= 12'b001000011001;
		12'd3585:BCD_Out <= 12'b001000011001;
		12'd3586:BCD_Out <= 12'b001000011001;
		12'd3587:BCD_Out <= 12'b001000011001;
		12'd3588:BCD_Out <= 12'b001000011001;
		12'd3589:BCD_Out <= 12'b001000011001;
		12'd3590:BCD_Out <= 12'b001000011001;
		12'd3591:BCD_Out <= 12'b001000011001;
		12'd3592:BCD_Out <= 12'b001000011001;
		12'd3593:BCD_Out <= 12'b001000011001;
		12'd3594:BCD_Out <= 12'b001000011001;
		12'd3595:BCD_Out <= 12'b001000011001;
		12'd3596:BCD_Out <= 12'b001000100000;
		12'd3597:BCD_Out <= 12'b001000100000;
		12'd3598:BCD_Out <= 12'b001000100000;
		12'd3599:BCD_Out <= 12'b001000100000;
		12'd3600:BCD_Out <= 12'b001000100000;
		12'd3601:BCD_Out <= 12'b001000100000;
		12'd3602:BCD_Out <= 12'b001000100000;
		12'd3603:BCD_Out <= 12'b001000100000;
		12'd3604:BCD_Out <= 12'b001000100000;
		12'd3605:BCD_Out <= 12'b001000100000;
		12'd3606:BCD_Out <= 12'b001000100000;
		12'd3607:BCD_Out <= 12'b001000100000;
		12'd3608:BCD_Out <= 12'b001000100000;
		12'd3609:BCD_Out <= 12'b001000100000;
		12'd3610:BCD_Out <= 12'b001000100000;
		12'd3611:BCD_Out <= 12'b001000100000;
		12'd3612:BCD_Out <= 12'b001000100001;
		12'd3613:BCD_Out <= 12'b001000100001;
		12'd3614:BCD_Out <= 12'b001000100001;
		12'd3615:BCD_Out <= 12'b001000100001;
		12'd3616:BCD_Out <= 12'b001000100001;
		12'd3617:BCD_Out <= 12'b001000100001;
		12'd3618:BCD_Out <= 12'b001000100001;
		12'd3619:BCD_Out <= 12'b001000100001;
		12'd3620:BCD_Out <= 12'b001000100001;
		12'd3621:BCD_Out <= 12'b001000100001;
		12'd3622:BCD_Out <= 12'b001000100001;
		12'd3623:BCD_Out <= 12'b001000100001;
		12'd3624:BCD_Out <= 12'b001000100001;
		12'd3625:BCD_Out <= 12'b001000100001;
		12'd3626:BCD_Out <= 12'b001000100001;
		12'd3627:BCD_Out <= 12'b001000100001;
		12'd3628:BCD_Out <= 12'b001000100001;
		12'd3629:BCD_Out <= 12'b001000100010;
		12'd3630:BCD_Out <= 12'b001000100010;
		12'd3631:BCD_Out <= 12'b001000100010;
		12'd3632:BCD_Out <= 12'b001000100010;
		12'd3633:BCD_Out <= 12'b001000100010;
		12'd3634:BCD_Out <= 12'b001000100010;
		12'd3635:BCD_Out <= 12'b001000100010;
		12'd3636:BCD_Out <= 12'b001000100010;
		12'd3637:BCD_Out <= 12'b001000100010;
		12'd3638:BCD_Out <= 12'b001000100010;
		12'd3639:BCD_Out <= 12'b001000100010;
		12'd3640:BCD_Out <= 12'b001000100010;
		12'd3641:BCD_Out <= 12'b001000100010;
		12'd3642:BCD_Out <= 12'b001000100010;
		12'd3643:BCD_Out <= 12'b001000100010;
		12'd3644:BCD_Out <= 12'b001000100010;
		12'd3645:BCD_Out <= 12'b001000100011;
		12'd3646:BCD_Out <= 12'b001000100011;
		12'd3647:BCD_Out <= 12'b001000100011;
		12'd3648:BCD_Out <= 12'b001000100011;
		12'd3649:BCD_Out <= 12'b001000100011;
		12'd3650:BCD_Out <= 12'b001000100011;
		12'd3651:BCD_Out <= 12'b001000100011;
		12'd3652:BCD_Out <= 12'b001000100011;
		12'd3653:BCD_Out <= 12'b001000100011;
		12'd3654:BCD_Out <= 12'b001000100011;
		12'd3655:BCD_Out <= 12'b001000100011;
		12'd3656:BCD_Out <= 12'b001000100011;
		12'd3657:BCD_Out <= 12'b001000100011;
		12'd3658:BCD_Out <= 12'b001000100011;
		12'd3659:BCD_Out <= 12'b001000100011;
		12'd3660:BCD_Out <= 12'b001000100011;
		12'd3661:BCD_Out <= 12'b001000100100;
		12'd3662:BCD_Out <= 12'b001000100100;
		12'd3663:BCD_Out <= 12'b001000100100;
		12'd3664:BCD_Out <= 12'b001000100100;
		12'd3665:BCD_Out <= 12'b001000100100;
		12'd3666:BCD_Out <= 12'b001000100100;
		12'd3667:BCD_Out <= 12'b001000100100;
		12'd3668:BCD_Out <= 12'b001000100100;
		12'd3669:BCD_Out <= 12'b001000100100;
		12'd3670:BCD_Out <= 12'b001000100100;
		12'd3671:BCD_Out <= 12'b001000100100;
		12'd3672:BCD_Out <= 12'b001000100100;
		12'd3673:BCD_Out <= 12'b001000100100;
		12'd3674:BCD_Out <= 12'b001000100100;
		12'd3675:BCD_Out <= 12'b001000100100;
		12'd3676:BCD_Out <= 12'b001000100100;
		12'd3677:BCD_Out <= 12'b001000100100;
		12'd3678:BCD_Out <= 12'b001000100101;
		12'd3679:BCD_Out <= 12'b001000100101;
		12'd3680:BCD_Out <= 12'b001000100101;
		12'd3681:BCD_Out <= 12'b001000100101;
		12'd3682:BCD_Out <= 12'b001000100101;
		12'd3683:BCD_Out <= 12'b001000100101;
		12'd3684:BCD_Out <= 12'b001000100101;
		12'd3685:BCD_Out <= 12'b001000100101;
		12'd3686:BCD_Out <= 12'b001000100101;
		12'd3687:BCD_Out <= 12'b001000100101;
		12'd3688:BCD_Out <= 12'b001000100101;
		12'd3689:BCD_Out <= 12'b001000100101;
		12'd3690:BCD_Out <= 12'b001000100101;
		12'd3691:BCD_Out <= 12'b001000100101;
		12'd3692:BCD_Out <= 12'b001000100101;
		12'd3693:BCD_Out <= 12'b001000100101;
		12'd3694:BCD_Out <= 12'b001000100110;
		12'd3695:BCD_Out <= 12'b001000100110;
		12'd3696:BCD_Out <= 12'b001000100110;
		12'd3697:BCD_Out <= 12'b001000100110;
		12'd3698:BCD_Out <= 12'b001000100110;
		12'd3699:BCD_Out <= 12'b001000100110;
		12'd3700:BCD_Out <= 12'b001000100110;
		12'd3701:BCD_Out <= 12'b001000100110;
		12'd3702:BCD_Out <= 12'b001000100110;
		12'd3703:BCD_Out <= 12'b001000100110;
		12'd3704:BCD_Out <= 12'b001000100110;
		12'd3705:BCD_Out <= 12'b001000100110;
		12'd3706:BCD_Out <= 12'b001000100110;
		12'd3707:BCD_Out <= 12'b001000100110;
		12'd3708:BCD_Out <= 12'b001000100110;
		12'd3709:BCD_Out <= 12'b001000100110;
		12'd3710:BCD_Out <= 12'b001000100110;
		12'd3711:BCD_Out <= 12'b001000100111;
		12'd3712:BCD_Out <= 12'b001000100111;
		12'd3713:BCD_Out <= 12'b001000100111;
		12'd3714:BCD_Out <= 12'b001000100111;
		12'd3715:BCD_Out <= 12'b001000100111;
		12'd3716:BCD_Out <= 12'b001000100111;
		12'd3717:BCD_Out <= 12'b001000100111;
		12'd3718:BCD_Out <= 12'b001000100111;
		12'd3719:BCD_Out <= 12'b001000100111;
		12'd3720:BCD_Out <= 12'b001000100111;
		12'd3721:BCD_Out <= 12'b001000100111;
		12'd3722:BCD_Out <= 12'b001000100111;
		12'd3723:BCD_Out <= 12'b001000100111;
		12'd3724:BCD_Out <= 12'b001000100111;
		12'd3725:BCD_Out <= 12'b001000100111;
		12'd3726:BCD_Out <= 12'b001000100111;
		12'd3727:BCD_Out <= 12'b001000101000;
		12'd3728:BCD_Out <= 12'b001000101000;
		12'd3729:BCD_Out <= 12'b001000101000;
		12'd3730:BCD_Out <= 12'b001000101000;
		12'd3731:BCD_Out <= 12'b001000101000;
		12'd3732:BCD_Out <= 12'b001000101000;
		12'd3733:BCD_Out <= 12'b001000101000;
		12'd3734:BCD_Out <= 12'b001000101000;
		12'd3735:BCD_Out <= 12'b001000101000;
		12'd3736:BCD_Out <= 12'b001000101000;
		12'd3737:BCD_Out <= 12'b001000101000;
		12'd3738:BCD_Out <= 12'b001000101000;
		12'd3739:BCD_Out <= 12'b001000101000;
		12'd3740:BCD_Out <= 12'b001000101000;
		12'd3741:BCD_Out <= 12'b001000101000;
		12'd3742:BCD_Out <= 12'b001000101000;
		12'd3743:BCD_Out <= 12'b001000101001;
		12'd3744:BCD_Out <= 12'b001000101001;
		12'd3745:BCD_Out <= 12'b001000101001;
		12'd3746:BCD_Out <= 12'b001000101001;
		12'd3747:BCD_Out <= 12'b001000101001;
		12'd3748:BCD_Out <= 12'b001000101001;
		12'd3749:BCD_Out <= 12'b001000101001;
		12'd3750:BCD_Out <= 12'b001000101001;
		12'd3751:BCD_Out <= 12'b001000101001;
		12'd3752:BCD_Out <= 12'b001000101001;
		12'd3753:BCD_Out <= 12'b001000101001;
		12'd3754:BCD_Out <= 12'b001000101001;
		12'd3755:BCD_Out <= 12'b001000101001;
		12'd3756:BCD_Out <= 12'b001000101001;
		12'd3757:BCD_Out <= 12'b001000101001;
		12'd3758:BCD_Out <= 12'b001000101001;
		12'd3759:BCD_Out <= 12'b001000101001;
		12'd3760:BCD_Out <= 12'b001000110000;
		12'd3761:BCD_Out <= 12'b001000110000;
		12'd3762:BCD_Out <= 12'b001000110000;
		12'd3763:BCD_Out <= 12'b001000110000;
		12'd3764:BCD_Out <= 12'b001000110000;
		12'd3765:BCD_Out <= 12'b001000110000;
		12'd3766:BCD_Out <= 12'b001000110000;
		12'd3767:BCD_Out <= 12'b001000110000;
		12'd3768:BCD_Out <= 12'b001000110000;
		12'd3769:BCD_Out <= 12'b001000110000;
		12'd3770:BCD_Out <= 12'b001000110000;
		12'd3771:BCD_Out <= 12'b001000110000;
		12'd3772:BCD_Out <= 12'b001000110000;
		12'd3773:BCD_Out <= 12'b001000110000;
		12'd3774:BCD_Out <= 12'b001000110000;
		12'd3775:BCD_Out <= 12'b001000110000;
		12'd3776:BCD_Out <= 12'b001000110001;
		12'd3777:BCD_Out <= 12'b001000110001;
		12'd3778:BCD_Out <= 12'b001000110001;
		12'd3779:BCD_Out <= 12'b001000110001;
		12'd3780:BCD_Out <= 12'b001000110001;
		12'd3781:BCD_Out <= 12'b001000110001;
		12'd3782:BCD_Out <= 12'b001000110001;
		12'd3783:BCD_Out <= 12'b001000110001;
		12'd3784:BCD_Out <= 12'b001000110001;
		12'd3785:BCD_Out <= 12'b001000110001;
		12'd3786:BCD_Out <= 12'b001000110001;
		12'd3787:BCD_Out <= 12'b001000110001;
		12'd3788:BCD_Out <= 12'b001000110001;
		12'd3789:BCD_Out <= 12'b001000110001;
		12'd3790:BCD_Out <= 12'b001000110001;
		12'd3791:BCD_Out <= 12'b001000110001;
		12'd3792:BCD_Out <= 12'b001000110010;
		12'd3793:BCD_Out <= 12'b001000110010;
		12'd3794:BCD_Out <= 12'b001000110010;
		12'd3795:BCD_Out <= 12'b001000110010;
		12'd3796:BCD_Out <= 12'b001000110010;
		12'd3797:BCD_Out <= 12'b001000110010;
		12'd3798:BCD_Out <= 12'b001000110010;
		12'd3799:BCD_Out <= 12'b001000110010;
		12'd3800:BCD_Out <= 12'b001000110010;
		12'd3801:BCD_Out <= 12'b001000110010;
		12'd3802:BCD_Out <= 12'b001000110010;
		12'd3803:BCD_Out <= 12'b001000110010;
		12'd3804:BCD_Out <= 12'b001000110010;
		12'd3805:BCD_Out <= 12'b001000110010;
		12'd3806:BCD_Out <= 12'b001000110010;
		12'd3807:BCD_Out <= 12'b001000110010;
		12'd3808:BCD_Out <= 12'b001000110010;
		12'd3809:BCD_Out <= 12'b001000110011;
		12'd3810:BCD_Out <= 12'b001000110011;
		12'd3811:BCD_Out <= 12'b001000110011;
		12'd3812:BCD_Out <= 12'b001000110011;
		12'd3813:BCD_Out <= 12'b001000110011;
		12'd3814:BCD_Out <= 12'b001000110011;
		12'd3815:BCD_Out <= 12'b001000110011;
		12'd3816:BCD_Out <= 12'b001000110011;
		12'd3817:BCD_Out <= 12'b001000110011;
		12'd3818:BCD_Out <= 12'b001000110011;
		12'd3819:BCD_Out <= 12'b001000110011;
		12'd3820:BCD_Out <= 12'b001000110011;
		12'd3821:BCD_Out <= 12'b001000110011;
		12'd3822:BCD_Out <= 12'b001000110011;
		12'd3823:BCD_Out <= 12'b001000110011;
		12'd3824:BCD_Out <= 12'b001000110011;
		12'd3825:BCD_Out <= 12'b001000110100;
		12'd3826:BCD_Out <= 12'b001000110100;
		12'd3827:BCD_Out <= 12'b001000110100;
		12'd3828:BCD_Out <= 12'b001000110100;
		12'd3829:BCD_Out <= 12'b001000110100;
		12'd3830:BCD_Out <= 12'b001000110100;
		12'd3831:BCD_Out <= 12'b001000110100;
		12'd3832:BCD_Out <= 12'b001000110100;
		12'd3833:BCD_Out <= 12'b001000110100;
		12'd3834:BCD_Out <= 12'b001000110100;
		12'd3835:BCD_Out <= 12'b001000110100;
		12'd3836:BCD_Out <= 12'b001000110100;
		12'd3837:BCD_Out <= 12'b001000110100;
		12'd3838:BCD_Out <= 12'b001000110100;
		12'd3839:BCD_Out <= 12'b001000110100;
		12'd3840:BCD_Out <= 12'b001000110100;
		12'd3841:BCD_Out <= 12'b001000110100;
		12'd3842:BCD_Out <= 12'b001000110101;
		12'd3843:BCD_Out <= 12'b001000110101;
		12'd3844:BCD_Out <= 12'b001000110101;
		12'd3845:BCD_Out <= 12'b001000110101;
		12'd3846:BCD_Out <= 12'b001000110101;
		12'd3847:BCD_Out <= 12'b001000110101;
		12'd3848:BCD_Out <= 12'b001000110101;
		12'd3849:BCD_Out <= 12'b001000110101;
		12'd3850:BCD_Out <= 12'b001000110101;
		12'd3851:BCD_Out <= 12'b001000110101;
		12'd3852:BCD_Out <= 12'b001000110101;
		12'd3853:BCD_Out <= 12'b001000110101;
		12'd3854:BCD_Out <= 12'b001000110101;
		12'd3855:BCD_Out <= 12'b001000110101;
		12'd3856:BCD_Out <= 12'b001000110101;
		12'd3857:BCD_Out <= 12'b001000110101;
		12'd3858:BCD_Out <= 12'b001000110110;
		12'd3859:BCD_Out <= 12'b001000110110;
		12'd3860:BCD_Out <= 12'b001000110110;
		12'd3861:BCD_Out <= 12'b001000110110;
		12'd3862:BCD_Out <= 12'b001000110110;
		12'd3863:BCD_Out <= 12'b001000110110;
		12'd3864:BCD_Out <= 12'b001000110110;
		12'd3865:BCD_Out <= 12'b001000110110;
		12'd3866:BCD_Out <= 12'b001000110110;
		12'd3867:BCD_Out <= 12'b001000110110;
		12'd3868:BCD_Out <= 12'b001000110110;
		12'd3869:BCD_Out <= 12'b001000110110;
		12'd3870:BCD_Out <= 12'b001000110110;
		12'd3871:BCD_Out <= 12'b001000110110;
		12'd3872:BCD_Out <= 12'b001000110110;
		12'd3873:BCD_Out <= 12'b001000110110;
		12'd3874:BCD_Out <= 12'b001000110111;
		12'd3875:BCD_Out <= 12'b001000110111;
		12'd3876:BCD_Out <= 12'b001000110111;
		12'd3877:BCD_Out <= 12'b001000110111;
		12'd3878:BCD_Out <= 12'b001000110111;
		12'd3879:BCD_Out <= 12'b001000110111;
		12'd3880:BCD_Out <= 12'b001000110111;
		12'd3881:BCD_Out <= 12'b001000110111;
		12'd3882:BCD_Out <= 12'b001000110111;
		12'd3883:BCD_Out <= 12'b001000110111;
		12'd3884:BCD_Out <= 12'b001000110111;
		12'd3885:BCD_Out <= 12'b001000110111;
		12'd3886:BCD_Out <= 12'b001000110111;
		12'd3887:BCD_Out <= 12'b001000110111;
		12'd3888:BCD_Out <= 12'b001000110111;
		12'd3889:BCD_Out <= 12'b001000110111;
		12'd3890:BCD_Out <= 12'b001000110111;
		12'd3891:BCD_Out <= 12'b001000111000;
		12'd3892:BCD_Out <= 12'b001000111000;
		12'd3893:BCD_Out <= 12'b001000111000;
		12'd3894:BCD_Out <= 12'b001000111000;
		12'd3895:BCD_Out <= 12'b001000111000;
		12'd3896:BCD_Out <= 12'b001000111000;
		12'd3897:BCD_Out <= 12'b001000111000;
		12'd3898:BCD_Out <= 12'b001000111000;
		12'd3899:BCD_Out <= 12'b001000111000;
		12'd3900:BCD_Out <= 12'b001000111000;
		12'd3901:BCD_Out <= 12'b001000111000;
		12'd3902:BCD_Out <= 12'b001000111000;
		12'd3903:BCD_Out <= 12'b001000111000;
		12'd3904:BCD_Out <= 12'b001000111000;
		12'd3905:BCD_Out <= 12'b001000111000;
		12'd3906:BCD_Out <= 12'b001000111000;
		12'd3907:BCD_Out <= 12'b001000111001;
		12'd3908:BCD_Out <= 12'b001000111001;
		12'd3909:BCD_Out <= 12'b001000111001;
		12'd3910:BCD_Out <= 12'b001000111001;
		12'd3911:BCD_Out <= 12'b001000111001;
		12'd3912:BCD_Out <= 12'b001000111001;
		12'd3913:BCD_Out <= 12'b001000111001;
		12'd3914:BCD_Out <= 12'b001000111001;
		12'd3915:BCD_Out <= 12'b001000111001;
		12'd3916:BCD_Out <= 12'b001000111001;
		12'd3917:BCD_Out <= 12'b001000111001;
		12'd3918:BCD_Out <= 12'b001000111001;
		12'd3919:BCD_Out <= 12'b001000111001;
		12'd3920:BCD_Out <= 12'b001000111001;
		12'd3921:BCD_Out <= 12'b001000111001;
		12'd3922:BCD_Out <= 12'b001000111001;
		12'd3923:BCD_Out <= 12'b001000111001;
		12'd3924:BCD_Out <= 12'b001001000000;
		12'd3925:BCD_Out <= 12'b001001000000;
		12'd3926:BCD_Out <= 12'b001001000000;
		12'd3927:BCD_Out <= 12'b001001000000;
		12'd3928:BCD_Out <= 12'b001001000000;
		12'd3929:BCD_Out <= 12'b001001000000;
		12'd3930:BCD_Out <= 12'b001001000000;
		12'd3931:BCD_Out <= 12'b001001000000;
		12'd3932:BCD_Out <= 12'b001001000000;
		12'd3933:BCD_Out <= 12'b001001000000;
		12'd3934:BCD_Out <= 12'b001001000000;
		12'd3935:BCD_Out <= 12'b001001000000;
		12'd3936:BCD_Out <= 12'b001001000000;
		12'd3937:BCD_Out <= 12'b001001000000;
		12'd3938:BCD_Out <= 12'b001001000000;
		12'd3939:BCD_Out <= 12'b001001000000;
		12'd3940:BCD_Out <= 12'b001001000001;
		12'd3941:BCD_Out <= 12'b001001000001;
		12'd3942:BCD_Out <= 12'b001001000001;
		12'd3943:BCD_Out <= 12'b001001000001;
		12'd3944:BCD_Out <= 12'b001001000001;
		12'd3945:BCD_Out <= 12'b001001000001;
		12'd3946:BCD_Out <= 12'b001001000001;
		12'd3947:BCD_Out <= 12'b001001000001;
		12'd3948:BCD_Out <= 12'b001001000001;
		12'd3949:BCD_Out <= 12'b001001000001;
		12'd3950:BCD_Out <= 12'b001001000001;
		12'd3951:BCD_Out <= 12'b001001000001;
		12'd3952:BCD_Out <= 12'b001001000001;
		12'd3953:BCD_Out <= 12'b001001000001;
		12'd3954:BCD_Out <= 12'b001001000001;
		12'd3955:BCD_Out <= 12'b001001000001;
		12'd3956:BCD_Out <= 12'b001001000010;
		12'd3957:BCD_Out <= 12'b001001000010;
		12'd3958:BCD_Out <= 12'b001001000010;
		12'd3959:BCD_Out <= 12'b001001000010;
		12'd3960:BCD_Out <= 12'b001001000010;
		12'd3961:BCD_Out <= 12'b001001000010;
		12'd3962:BCD_Out <= 12'b001001000010;
		12'd3963:BCD_Out <= 12'b001001000010;
		12'd3964:BCD_Out <= 12'b001001000010;
		12'd3965:BCD_Out <= 12'b001001000010;
		12'd3966:BCD_Out <= 12'b001001000010;
		12'd3967:BCD_Out <= 12'b001001000010;
		12'd3968:BCD_Out <= 12'b001001000010;
		12'd3969:BCD_Out <= 12'b001001000010;
		12'd3970:BCD_Out <= 12'b001001000010;
		12'd3971:BCD_Out <= 12'b001001000010;
		12'd3972:BCD_Out <= 12'b001001000010;
		12'd3973:BCD_Out <= 12'b001001000011;
		12'd3974:BCD_Out <= 12'b001001000011;
		12'd3975:BCD_Out <= 12'b001001000011;
		12'd3976:BCD_Out <= 12'b001001000011;
		12'd3977:BCD_Out <= 12'b001001000011;
		12'd3978:BCD_Out <= 12'b001001000011;
		12'd3979:BCD_Out <= 12'b001001000011;
		12'd3980:BCD_Out <= 12'b001001000011;
		12'd3981:BCD_Out <= 12'b001001000011;
		12'd3982:BCD_Out <= 12'b001001000011;
		12'd3983:BCD_Out <= 12'b001001000011;
		12'd3984:BCD_Out <= 12'b001001000011;
		12'd3985:BCD_Out <= 12'b001001000011;
		12'd3986:BCD_Out <= 12'b001001000011;
		12'd3987:BCD_Out <= 12'b001001000011;
		12'd3988:BCD_Out <= 12'b001001000011;
		12'd3989:BCD_Out <= 12'b001001000100;
		12'd3990:BCD_Out <= 12'b001001000100;
		12'd3991:BCD_Out <= 12'b001001000100;
		12'd3992:BCD_Out <= 12'b001001000100;
		12'd3993:BCD_Out <= 12'b001001000100;
		12'd3994:BCD_Out <= 12'b001001000100;
		12'd3995:BCD_Out <= 12'b001001000100;
		12'd3996:BCD_Out <= 12'b001001000100;
		12'd3997:BCD_Out <= 12'b001001000100;
		12'd3998:BCD_Out <= 12'b001001000100;
		12'd3999:BCD_Out <= 12'b001001000100;
		12'd4000:BCD_Out <= 12'b001001000100;
		12'd4001:BCD_Out <= 12'b001001000100;
		12'd4002:BCD_Out <= 12'b001001000100;
		12'd4003:BCD_Out <= 12'b001001000100;
		12'd4004:BCD_Out <= 12'b001001000100;
		12'd4005:BCD_Out <= 12'b001001000101;
		12'd4006:BCD_Out <= 12'b001001000101;
		12'd4007:BCD_Out <= 12'b001001000101;
		12'd4008:BCD_Out <= 12'b001001000101;
		12'd4009:BCD_Out <= 12'b001001000101;
		12'd4010:BCD_Out <= 12'b001001000101;
		12'd4011:BCD_Out <= 12'b001001000101;
		12'd4012:BCD_Out <= 12'b001001000101;
		12'd4013:BCD_Out <= 12'b001001000101;
		12'd4014:BCD_Out <= 12'b001001000101;
		12'd4015:BCD_Out <= 12'b001001000101;
		12'd4016:BCD_Out <= 12'b001001000101;
		12'd4017:BCD_Out <= 12'b001001000101;
		12'd4018:BCD_Out <= 12'b001001000101;
		12'd4019:BCD_Out <= 12'b001001000101;
		12'd4020:BCD_Out <= 12'b001001000101;
		12'd4021:BCD_Out <= 12'b001001000101;
		12'd4022:BCD_Out <= 12'b001001000110;
		12'd4023:BCD_Out <= 12'b001001000110;
		12'd4024:BCD_Out <= 12'b001001000110;
		12'd4025:BCD_Out <= 12'b001001000110;
		12'd4026:BCD_Out <= 12'b001001000110;
		12'd4027:BCD_Out <= 12'b001001000110;
		12'd4028:BCD_Out <= 12'b001001000110;
		12'd4029:BCD_Out <= 12'b001001000110;
		12'd4030:BCD_Out <= 12'b001001000110;
		12'd4031:BCD_Out <= 12'b001001000110;
		12'd4032:BCD_Out <= 12'b001001000110;
		12'd4033:BCD_Out <= 12'b001001000110;
		12'd4034:BCD_Out <= 12'b001001000110;
		12'd4035:BCD_Out <= 12'b001001000110;
		12'd4036:BCD_Out <= 12'b001001000110;
		12'd4037:BCD_Out <= 12'b001001000110;
		12'd4038:BCD_Out <= 12'b001001000111;
		12'd4039:BCD_Out <= 12'b001001000111;
		12'd4040:BCD_Out <= 12'b001001000111;
		12'd4041:BCD_Out <= 12'b001001000111;
		12'd4042:BCD_Out <= 12'b001001000111;
		12'd4043:BCD_Out <= 12'b001001000111;
		12'd4044:BCD_Out <= 12'b001001000111;
		12'd4045:BCD_Out <= 12'b001001000111;
		12'd4046:BCD_Out <= 12'b001001000111;
		12'd4047:BCD_Out <= 12'b001001000111;
		12'd4048:BCD_Out <= 12'b001001000111;
		12'd4049:BCD_Out <= 12'b001001000111;
		12'd4050:BCD_Out <= 12'b001001000111;
		12'd4051:BCD_Out <= 12'b001001000111;
		12'd4052:BCD_Out <= 12'b001001000111;
		12'd4053:BCD_Out <= 12'b001001000111;
		12'd4054:BCD_Out <= 12'b001001000111;
		12'd4055:BCD_Out <= 12'b001001001000;
		12'd4056:BCD_Out <= 12'b001001001000;
		12'd4057:BCD_Out <= 12'b001001001000;
		12'd4058:BCD_Out <= 12'b001001001000;
		12'd4059:BCD_Out <= 12'b001001001000;
		12'd4060:BCD_Out <= 12'b001001001000;
		12'd4061:BCD_Out <= 12'b001001001000;
		12'd4062:BCD_Out <= 12'b001001001000;
		12'd4063:BCD_Out <= 12'b001001001000;
		12'd4064:BCD_Out <= 12'b001001001000;
		12'd4065:BCD_Out <= 12'b001001001000;
		12'd4066:BCD_Out <= 12'b001001001000;
		12'd4067:BCD_Out <= 12'b001001001000;
		12'd4068:BCD_Out <= 12'b001001001000;
		12'd4069:BCD_Out <= 12'b001001001000;
		12'd4070:BCD_Out <= 12'b001001001000;
		12'd4071:BCD_Out <= 12'b001001001001;
		12'd4072:BCD_Out <= 12'b001001001001;
		12'd4073:BCD_Out <= 12'b001001001001;
		12'd4074:BCD_Out <= 12'b001001001001;
		12'd4075:BCD_Out <= 12'b001001001001;
		12'd4076:BCD_Out <= 12'b001001001001;
		12'd4077:BCD_Out <= 12'b001001001001;
		12'd4078:BCD_Out <= 12'b001001001001;
		12'd4079:BCD_Out <= 12'b001001001001;
		12'd4080:BCD_Out <= 12'b001001001001;
		12'd4081:BCD_Out <= 12'b001001001001;
		12'd4082:BCD_Out <= 12'b001001001001;
		12'd4083:BCD_Out <= 12'b001001001001;
		12'd4084:BCD_Out <= 12'b001001001001;
		12'd4085:BCD_Out <= 12'b001001001001;
		12'd4086:BCD_Out <= 12'b001001001001;
		12'd4087:BCD_Out <= 12'b001001010000;
		12'd4088:BCD_Out <= 12'b001001010000;
		12'd4089:BCD_Out <= 12'b001001010000;
		12'd4090:BCD_Out <= 12'b001001010000;
		12'd4091:BCD_Out <= 12'b001001010000;
		12'd4092:BCD_Out <= 12'b001001010000;
		12'd4093:BCD_Out <= 12'b001001010000;
		12'd4094:BCD_Out <= 12'b001001010000;
		12'd4095:BCD_Out <= 12'b001001010000;
		default:BCD_Out <= 12'b000000000000;
	endcase
end

endmodule
